magic
tech scmos
timestamp 1731962781
<< nwell >>
rect 1772 384 1826 446
rect 1834 314 1861 376
rect 2150 307 2202 334
rect 2248 302 2275 347
rect 2150 256 2202 283
rect 2402 189 2429 285
rect 2451 192 2478 237
rect -3142 -2166 -3090 -2139
rect -3044 -2171 -3017 -2126
rect -3142 -2217 -3090 -2190
rect -2940 -2213 -2886 -2151
rect -2878 -2283 -2851 -2221
rect -2795 -2251 -2741 -2189
rect -3158 -2374 -3104 -2312
rect -2733 -2321 -2706 -2259
rect -2602 -2267 -2548 -2205
rect -2456 -2265 -2402 -2203
rect -2312 -2269 -2258 -2207
rect -2157 -2271 -2103 -2209
rect -2540 -2337 -2513 -2275
rect -2394 -2335 -2367 -2273
rect -2250 -2339 -2223 -2277
rect -2022 -2279 -1968 -2217
rect -2095 -2341 -2068 -2279
rect -1960 -2349 -1933 -2287
rect -1861 -2369 -1834 -2273
rect -1812 -2366 -1785 -2321
rect -3096 -2444 -3069 -2382
rect -1699 -2425 -1672 -2329
rect -1650 -2422 -1623 -2377
rect -1541 -2481 -1514 -2385
rect -1492 -2478 -1465 -2433
rect -1375 -2557 -1348 -2461
rect -1326 -2554 -1299 -2509
rect -3136 -3017 -3084 -2990
rect -3038 -3022 -3011 -2977
rect -2932 -3028 -2878 -2966
rect -2763 -3027 -2709 -2965
rect -2599 -3025 -2545 -2963
rect -2459 -3027 -2405 -2965
rect -3136 -3068 -3084 -3041
rect -2870 -3098 -2843 -3036
rect -2701 -3097 -2674 -3035
rect -2537 -3095 -2510 -3033
rect -2397 -3097 -2370 -3035
rect -2308 -3040 -2254 -2978
rect -2246 -3110 -2219 -3048
rect -1998 -3116 -1971 -3020
rect -1949 -3113 -1922 -3068
rect -3165 -3289 -3111 -3227
rect -2145 -3244 -2091 -3182
rect -3103 -3359 -3076 -3297
rect -2083 -3314 -2056 -3252
rect -1864 -3326 -1837 -3230
rect -1815 -3323 -1788 -3278
rect -1717 -3486 -1690 -3390
rect -1668 -3483 -1641 -3438
rect -1505 -3450 -1481 -3418
rect -1505 -3505 -1463 -3473
rect -3136 -3785 -3084 -3758
rect -3038 -3790 -3011 -3745
rect -2911 -3801 -2857 -3739
rect -3136 -3836 -3084 -3809
rect -2849 -3871 -2822 -3809
rect -2910 -4006 -2856 -3944
rect -2745 -3976 -2718 -3880
rect -2696 -3973 -2669 -3928
rect -2848 -4076 -2821 -4014
rect -3171 -4138 -3117 -4076
rect -2599 -4089 -2572 -3993
rect -2550 -4086 -2523 -4041
rect -2423 -4061 -2399 -4029
rect -2423 -4116 -2381 -4084
rect -3109 -4208 -3082 -4146
rect 702 -4161 726 -4129
rect 702 -4216 744 -4184
rect -3158 -4547 -3106 -4520
rect -3060 -4552 -3033 -4507
rect -3158 -4598 -3106 -4571
rect -2999 -4581 -2945 -4519
rect -2937 -4651 -2910 -4589
rect -3168 -4761 -3114 -4699
rect -3106 -4831 -3079 -4769
rect -2851 -4819 -2824 -4723
rect -2802 -4816 -2775 -4771
rect -2615 -4785 -2591 -4753
rect -2615 -4840 -2573 -4808
rect -2943 -4901 -2919 -4869
rect -2943 -4956 -2901 -4924
<< ntransistor >>
rect 1804 318 1806 338
rect 2120 319 2130 321
rect 2225 307 2227 317
rect 1847 284 1849 295
rect 1804 263 1806 283
rect 2225 274 2227 284
rect 2261 282 2263 292
rect 2120 268 2130 270
rect 2464 172 2466 182
rect 2400 162 2402 172
rect 2433 162 2435 172
rect -3172 -2154 -3162 -2152
rect -3067 -2166 -3065 -2158
rect -3067 -2199 -3065 -2189
rect -3031 -2191 -3029 -2181
rect -3172 -2205 -3162 -2203
rect -2908 -2279 -2906 -2259
rect -2865 -2313 -2863 -2302
rect -2908 -2334 -2906 -2314
rect -2763 -2317 -2761 -2297
rect -2570 -2333 -2568 -2313
rect -2720 -2351 -2718 -2340
rect -2763 -2372 -2761 -2352
rect -2424 -2331 -2422 -2311
rect -2280 -2335 -2278 -2315
rect -2527 -2367 -2525 -2356
rect -2381 -2365 -2379 -2354
rect -2125 -2337 -2123 -2317
rect -2570 -2388 -2568 -2368
rect -2424 -2386 -2422 -2366
rect -2237 -2369 -2235 -2358
rect -1990 -2345 -1988 -2325
rect -2280 -2390 -2278 -2370
rect -2082 -2371 -2080 -2360
rect -2125 -2392 -2123 -2372
rect -1947 -2379 -1945 -2368
rect -3126 -2440 -3124 -2420
rect -1990 -2400 -1988 -2380
rect -1799 -2386 -1797 -2376
rect -1863 -2396 -1861 -2386
rect -1830 -2396 -1828 -2386
rect -1637 -2442 -1635 -2432
rect -1701 -2452 -1699 -2442
rect -1668 -2452 -1666 -2442
rect -3083 -2474 -3081 -2463
rect -3126 -2495 -3124 -2475
rect -1479 -2498 -1477 -2488
rect -1543 -2508 -1541 -2498
rect -1510 -2508 -1508 -2498
rect -1313 -2574 -1311 -2564
rect -1377 -2584 -1375 -2574
rect -1344 -2584 -1342 -2574
rect -3166 -3005 -3156 -3003
rect -3061 -3017 -3059 -3009
rect -3061 -3050 -3059 -3040
rect -3025 -3042 -3023 -3032
rect -3166 -3056 -3156 -3054
rect -2900 -3094 -2898 -3074
rect -2731 -3093 -2729 -3073
rect -2567 -3091 -2565 -3071
rect -2427 -3093 -2425 -3073
rect -2857 -3128 -2855 -3117
rect -2688 -3127 -2686 -3116
rect -2524 -3125 -2522 -3114
rect -2276 -3106 -2274 -3086
rect -2900 -3149 -2898 -3129
rect -2731 -3148 -2729 -3128
rect -2567 -3146 -2565 -3126
rect -2384 -3127 -2382 -3116
rect -2427 -3148 -2425 -3128
rect -2233 -3140 -2231 -3129
rect -1936 -3133 -1934 -3123
rect -2276 -3161 -2274 -3141
rect -2000 -3143 -1998 -3133
rect -1967 -3143 -1965 -3133
rect -2113 -3310 -2111 -3290
rect -3133 -3355 -3131 -3335
rect -2070 -3344 -2068 -3333
rect -1802 -3343 -1800 -3333
rect -2113 -3365 -2111 -3345
rect -1866 -3353 -1864 -3343
rect -1833 -3353 -1831 -3343
rect -3090 -3389 -3088 -3378
rect -3133 -3410 -3131 -3390
rect -1494 -3467 -1492 -3457
rect -1655 -3503 -1653 -3493
rect -1719 -3513 -1717 -3503
rect -1686 -3513 -1684 -3503
rect -1494 -3521 -1492 -3511
rect -1476 -3521 -1474 -3511
rect -3166 -3773 -3156 -3771
rect -3061 -3785 -3059 -3777
rect -3061 -3818 -3059 -3808
rect -3025 -3810 -3023 -3800
rect -3166 -3824 -3156 -3822
rect -2879 -3867 -2877 -3847
rect -2836 -3901 -2834 -3890
rect -2879 -3922 -2877 -3902
rect -2683 -3993 -2681 -3983
rect -2747 -4003 -2745 -3993
rect -2714 -4003 -2712 -3993
rect -2878 -4072 -2876 -4052
rect -2835 -4106 -2833 -4095
rect -2412 -4078 -2410 -4068
rect -2537 -4106 -2535 -4096
rect -2878 -4127 -2876 -4107
rect -2601 -4116 -2599 -4106
rect -2568 -4116 -2566 -4106
rect -2412 -4132 -2410 -4122
rect -2394 -4132 -2392 -4122
rect -3139 -4204 -3137 -4184
rect 713 -4178 715 -4168
rect -3096 -4238 -3094 -4227
rect 713 -4232 715 -4222
rect 731 -4232 733 -4222
rect -3139 -4259 -3137 -4239
rect -3188 -4535 -3178 -4533
rect -3083 -4547 -3081 -4539
rect -3083 -4580 -3081 -4570
rect -3047 -4572 -3045 -4562
rect -3188 -4586 -3178 -4584
rect -2967 -4647 -2965 -4627
rect -2924 -4681 -2922 -4670
rect -2967 -4702 -2965 -4682
rect -3136 -4827 -3134 -4807
rect -2604 -4802 -2602 -4792
rect -2789 -4836 -2787 -4826
rect -2853 -4846 -2851 -4836
rect -2820 -4846 -2818 -4836
rect -3093 -4861 -3091 -4850
rect -2604 -4856 -2602 -4846
rect -2586 -4856 -2584 -4846
rect -3136 -4882 -3134 -4862
rect -2932 -4918 -2930 -4908
rect -2932 -4972 -2930 -4962
rect -2914 -4972 -2912 -4962
<< ptransistor >>
rect 1785 392 1787 412
rect 1812 392 1814 412
rect 1847 322 1849 362
rect 2158 319 2178 321
rect 2261 310 2263 330
rect 2158 268 2178 270
rect 2415 244 2417 264
rect 2415 197 2417 216
rect 2464 200 2466 220
rect -3134 -2154 -3114 -2152
rect -3031 -2163 -3029 -2143
rect -3134 -2205 -3114 -2203
rect -2927 -2205 -2925 -2185
rect -2900 -2205 -2898 -2185
rect -2865 -2275 -2863 -2235
rect -2782 -2243 -2780 -2223
rect -2755 -2243 -2753 -2223
rect -2589 -2259 -2587 -2239
rect -2562 -2259 -2560 -2239
rect -2443 -2257 -2441 -2237
rect -2416 -2257 -2414 -2237
rect -2720 -2313 -2718 -2273
rect -2299 -2261 -2297 -2241
rect -2272 -2261 -2270 -2241
rect -2527 -2329 -2525 -2289
rect -2144 -2263 -2142 -2243
rect -2117 -2263 -2115 -2243
rect -3145 -2366 -3143 -2346
rect -3118 -2366 -3116 -2346
rect -2381 -2327 -2379 -2287
rect -2009 -2271 -2007 -2251
rect -1982 -2271 -1980 -2251
rect -2237 -2331 -2235 -2291
rect -2082 -2333 -2080 -2293
rect -1947 -2341 -1945 -2301
rect -1848 -2314 -1846 -2294
rect -1848 -2361 -1846 -2342
rect -3083 -2436 -3081 -2396
rect -1799 -2358 -1797 -2338
rect -1686 -2370 -1684 -2350
rect -1686 -2417 -1684 -2398
rect -1637 -2414 -1635 -2394
rect -1528 -2426 -1526 -2406
rect -1528 -2473 -1526 -2454
rect -1479 -2470 -1477 -2450
rect -1362 -2502 -1360 -2482
rect -1362 -2549 -1360 -2530
rect -1313 -2546 -1311 -2526
rect -3128 -3005 -3108 -3003
rect -3025 -3014 -3023 -2994
rect -2919 -3020 -2917 -3000
rect -2892 -3020 -2890 -3000
rect -2750 -3019 -2748 -2999
rect -2723 -3019 -2721 -2999
rect -2586 -3017 -2584 -2997
rect -2559 -3017 -2557 -2997
rect -2446 -3019 -2444 -2999
rect -2419 -3019 -2417 -2999
rect -2295 -3032 -2293 -3012
rect -2268 -3032 -2266 -3012
rect -3128 -3056 -3108 -3054
rect -2857 -3090 -2855 -3050
rect -2688 -3089 -2686 -3049
rect -2524 -3087 -2522 -3047
rect -2384 -3089 -2382 -3049
rect -1985 -3061 -1983 -3041
rect -2233 -3102 -2231 -3062
rect -1985 -3108 -1983 -3089
rect -1936 -3105 -1934 -3085
rect -2132 -3236 -2130 -3216
rect -2105 -3236 -2103 -3216
rect -3152 -3281 -3150 -3261
rect -3125 -3281 -3123 -3261
rect -2070 -3306 -2068 -3266
rect -1851 -3271 -1849 -3251
rect -3090 -3351 -3088 -3311
rect -1851 -3318 -1849 -3299
rect -1802 -3315 -1800 -3295
rect -1704 -3431 -1702 -3411
rect -1704 -3478 -1702 -3459
rect -1494 -3444 -1492 -3424
rect -1655 -3475 -1653 -3455
rect -1494 -3499 -1492 -3479
rect -1476 -3499 -1474 -3479
rect -3128 -3773 -3108 -3771
rect -3025 -3782 -3023 -3762
rect -2898 -3793 -2896 -3773
rect -2871 -3793 -2869 -3773
rect -3128 -3824 -3108 -3822
rect -2836 -3863 -2834 -3823
rect -2732 -3921 -2730 -3901
rect -2732 -3968 -2730 -3949
rect -2897 -3998 -2895 -3978
rect -2870 -3998 -2868 -3978
rect -2683 -3965 -2681 -3945
rect -2835 -4068 -2833 -4028
rect -2586 -4034 -2584 -4014
rect -2586 -4081 -2584 -4062
rect -2412 -4055 -2410 -4035
rect -2537 -4078 -2535 -4058
rect -3158 -4130 -3156 -4110
rect -3131 -4130 -3129 -4110
rect -2412 -4110 -2410 -4090
rect -2394 -4110 -2392 -4090
rect 713 -4155 715 -4135
rect -3096 -4200 -3094 -4160
rect 713 -4210 715 -4190
rect 731 -4210 733 -4190
rect -3150 -4535 -3130 -4533
rect -3047 -4544 -3045 -4524
rect -2986 -4573 -2984 -4553
rect -2959 -4573 -2957 -4553
rect -3150 -4586 -3130 -4584
rect -2924 -4643 -2922 -4603
rect -3155 -4753 -3153 -4733
rect -3128 -4753 -3126 -4733
rect -2838 -4764 -2836 -4744
rect -3093 -4823 -3091 -4783
rect -2838 -4811 -2836 -4792
rect -2604 -4779 -2602 -4759
rect -2789 -4808 -2787 -4788
rect -2604 -4834 -2602 -4814
rect -2586 -4834 -2584 -4814
rect -2932 -4895 -2930 -4875
rect -2932 -4950 -2930 -4930
rect -2914 -4950 -2912 -4930
<< ndiffusion >>
rect 1803 318 1804 338
rect 1806 318 1807 338
rect 2120 321 2130 322
rect 2120 318 2130 319
rect 2224 307 2225 317
rect 2227 307 2228 317
rect 1846 284 1847 295
rect 1849 284 1850 295
rect 1803 263 1804 283
rect 1806 263 1807 283
rect 2120 270 2130 271
rect 2224 274 2225 284
rect 2227 274 2228 284
rect 2260 282 2261 292
rect 2263 282 2264 292
rect 2120 267 2130 268
rect 2463 172 2464 182
rect 2466 172 2467 182
rect 2399 162 2400 172
rect 2402 162 2403 172
rect 2432 162 2433 172
rect 2435 162 2436 172
rect -3172 -2152 -3162 -2151
rect -3172 -2155 -3162 -2154
rect -3068 -2166 -3067 -2158
rect -3065 -2166 -3064 -2158
rect -3172 -2203 -3162 -2202
rect -3068 -2199 -3067 -2189
rect -3065 -2199 -3064 -2189
rect -3032 -2191 -3031 -2181
rect -3029 -2191 -3028 -2181
rect -3172 -2206 -3162 -2205
rect -2909 -2279 -2908 -2259
rect -2906 -2279 -2905 -2259
rect -2866 -2313 -2865 -2302
rect -2863 -2313 -2862 -2302
rect -2909 -2334 -2908 -2314
rect -2906 -2334 -2905 -2314
rect -2764 -2317 -2763 -2297
rect -2761 -2317 -2760 -2297
rect -2571 -2333 -2570 -2313
rect -2568 -2333 -2567 -2313
rect -2721 -2351 -2720 -2340
rect -2718 -2351 -2717 -2340
rect -2764 -2372 -2763 -2352
rect -2761 -2372 -2760 -2352
rect -2425 -2331 -2424 -2311
rect -2422 -2331 -2421 -2311
rect -2281 -2335 -2280 -2315
rect -2278 -2335 -2277 -2315
rect -2528 -2367 -2527 -2356
rect -2525 -2367 -2524 -2356
rect -2382 -2365 -2381 -2354
rect -2379 -2365 -2378 -2354
rect -2126 -2337 -2125 -2317
rect -2123 -2337 -2122 -2317
rect -2571 -2388 -2570 -2368
rect -2568 -2388 -2567 -2368
rect -2425 -2386 -2424 -2366
rect -2422 -2386 -2421 -2366
rect -2238 -2369 -2237 -2358
rect -2235 -2369 -2234 -2358
rect -1991 -2345 -1990 -2325
rect -1988 -2345 -1987 -2325
rect -2281 -2390 -2280 -2370
rect -2278 -2390 -2277 -2370
rect -2083 -2371 -2082 -2360
rect -2080 -2371 -2079 -2360
rect -2126 -2392 -2125 -2372
rect -2123 -2392 -2122 -2372
rect -1948 -2379 -1947 -2368
rect -1945 -2379 -1944 -2368
rect -3127 -2440 -3126 -2420
rect -3124 -2440 -3123 -2420
rect -1991 -2400 -1990 -2380
rect -1988 -2400 -1987 -2380
rect -1800 -2386 -1799 -2376
rect -1797 -2386 -1796 -2376
rect -1864 -2396 -1863 -2386
rect -1861 -2396 -1860 -2386
rect -1831 -2396 -1830 -2386
rect -1828 -2396 -1827 -2386
rect -1638 -2442 -1637 -2432
rect -1635 -2442 -1634 -2432
rect -1702 -2452 -1701 -2442
rect -1699 -2452 -1698 -2442
rect -1669 -2452 -1668 -2442
rect -1666 -2452 -1665 -2442
rect -3084 -2474 -3083 -2463
rect -3081 -2474 -3080 -2463
rect -3127 -2495 -3126 -2475
rect -3124 -2495 -3123 -2475
rect -1480 -2498 -1479 -2488
rect -1477 -2498 -1476 -2488
rect -1544 -2508 -1543 -2498
rect -1541 -2508 -1540 -2498
rect -1511 -2508 -1510 -2498
rect -1508 -2508 -1507 -2498
rect -1314 -2574 -1313 -2564
rect -1311 -2574 -1310 -2564
rect -1378 -2584 -1377 -2574
rect -1375 -2584 -1374 -2574
rect -1345 -2584 -1344 -2574
rect -1342 -2584 -1341 -2574
rect -3166 -3003 -3156 -3002
rect -3166 -3006 -3156 -3005
rect -3062 -3017 -3061 -3009
rect -3059 -3017 -3058 -3009
rect -3166 -3054 -3156 -3053
rect -3062 -3050 -3061 -3040
rect -3059 -3050 -3058 -3040
rect -3026 -3042 -3025 -3032
rect -3023 -3042 -3022 -3032
rect -3166 -3057 -3156 -3056
rect -2901 -3094 -2900 -3074
rect -2898 -3094 -2897 -3074
rect -2732 -3093 -2731 -3073
rect -2729 -3093 -2728 -3073
rect -2568 -3091 -2567 -3071
rect -2565 -3091 -2564 -3071
rect -2428 -3093 -2427 -3073
rect -2425 -3093 -2424 -3073
rect -2858 -3128 -2857 -3117
rect -2855 -3128 -2854 -3117
rect -2689 -3127 -2688 -3116
rect -2686 -3127 -2685 -3116
rect -2525 -3125 -2524 -3114
rect -2522 -3125 -2521 -3114
rect -2277 -3106 -2276 -3086
rect -2274 -3106 -2273 -3086
rect -2901 -3149 -2900 -3129
rect -2898 -3149 -2897 -3129
rect -2732 -3148 -2731 -3128
rect -2729 -3148 -2728 -3128
rect -2568 -3146 -2567 -3126
rect -2565 -3146 -2564 -3126
rect -2385 -3127 -2384 -3116
rect -2382 -3127 -2381 -3116
rect -2428 -3148 -2427 -3128
rect -2425 -3148 -2424 -3128
rect -2234 -3140 -2233 -3129
rect -2231 -3140 -2230 -3129
rect -1937 -3133 -1936 -3123
rect -1934 -3133 -1933 -3123
rect -2277 -3161 -2276 -3141
rect -2274 -3161 -2273 -3141
rect -2001 -3143 -2000 -3133
rect -1998 -3143 -1997 -3133
rect -1968 -3143 -1967 -3133
rect -1965 -3143 -1964 -3133
rect -2114 -3310 -2113 -3290
rect -2111 -3310 -2110 -3290
rect -3134 -3355 -3133 -3335
rect -3131 -3355 -3130 -3335
rect -2071 -3344 -2070 -3333
rect -2068 -3344 -2067 -3333
rect -1803 -3343 -1802 -3333
rect -1800 -3343 -1799 -3333
rect -2114 -3365 -2113 -3345
rect -2111 -3365 -2110 -3345
rect -1867 -3353 -1866 -3343
rect -1864 -3353 -1863 -3343
rect -1834 -3353 -1833 -3343
rect -1831 -3353 -1830 -3343
rect -3091 -3389 -3090 -3378
rect -3088 -3389 -3087 -3378
rect -3134 -3410 -3133 -3390
rect -3131 -3410 -3130 -3390
rect -1499 -3463 -1494 -3457
rect -1495 -3467 -1494 -3463
rect -1492 -3461 -1491 -3457
rect -1492 -3467 -1487 -3461
rect -1656 -3503 -1655 -3493
rect -1653 -3503 -1652 -3493
rect -1720 -3513 -1719 -3503
rect -1717 -3513 -1716 -3503
rect -1687 -3513 -1686 -3503
rect -1684 -3513 -1683 -3503
rect -1499 -3517 -1494 -3511
rect -1495 -3521 -1494 -3517
rect -1492 -3515 -1491 -3511
rect -1492 -3521 -1487 -3515
rect -1477 -3515 -1476 -3511
rect -1481 -3521 -1476 -3515
rect -1474 -3515 -1473 -3511
rect -1474 -3521 -1469 -3515
rect -3166 -3771 -3156 -3770
rect -3166 -3774 -3156 -3773
rect -3062 -3785 -3061 -3777
rect -3059 -3785 -3058 -3777
rect -3166 -3822 -3156 -3821
rect -3062 -3818 -3061 -3808
rect -3059 -3818 -3058 -3808
rect -3026 -3810 -3025 -3800
rect -3023 -3810 -3022 -3800
rect -3166 -3825 -3156 -3824
rect -2880 -3867 -2879 -3847
rect -2877 -3867 -2876 -3847
rect -2837 -3901 -2836 -3890
rect -2834 -3901 -2833 -3890
rect -2880 -3922 -2879 -3902
rect -2877 -3922 -2876 -3902
rect -2684 -3993 -2683 -3983
rect -2681 -3993 -2680 -3983
rect -2748 -4003 -2747 -3993
rect -2745 -4003 -2744 -3993
rect -2715 -4003 -2714 -3993
rect -2712 -4003 -2711 -3993
rect -2879 -4072 -2878 -4052
rect -2876 -4072 -2875 -4052
rect -2836 -4106 -2835 -4095
rect -2833 -4106 -2832 -4095
rect -2417 -4074 -2412 -4068
rect -2413 -4078 -2412 -4074
rect -2410 -4072 -2409 -4068
rect -2410 -4078 -2405 -4072
rect -2538 -4106 -2537 -4096
rect -2535 -4106 -2534 -4096
rect -2879 -4127 -2878 -4107
rect -2876 -4127 -2875 -4107
rect -2602 -4116 -2601 -4106
rect -2599 -4116 -2598 -4106
rect -2569 -4116 -2568 -4106
rect -2566 -4116 -2565 -4106
rect -2417 -4128 -2412 -4122
rect -2413 -4132 -2412 -4128
rect -2410 -4126 -2409 -4122
rect -2410 -4132 -2405 -4126
rect -2395 -4126 -2394 -4122
rect -2399 -4132 -2394 -4126
rect -2392 -4126 -2391 -4122
rect -2392 -4132 -2387 -4126
rect -3140 -4204 -3139 -4184
rect -3137 -4204 -3136 -4184
rect 708 -4174 713 -4168
rect 712 -4178 713 -4174
rect 715 -4172 716 -4168
rect 715 -4178 720 -4172
rect -3097 -4238 -3096 -4227
rect -3094 -4238 -3093 -4227
rect 708 -4228 713 -4222
rect 712 -4232 713 -4228
rect 715 -4226 716 -4222
rect 715 -4232 720 -4226
rect 730 -4226 731 -4222
rect 726 -4232 731 -4226
rect 733 -4226 734 -4222
rect 733 -4232 738 -4226
rect -3140 -4259 -3139 -4239
rect -3137 -4259 -3136 -4239
rect -3188 -4533 -3178 -4532
rect -3188 -4536 -3178 -4535
rect -3084 -4547 -3083 -4539
rect -3081 -4547 -3080 -4539
rect -3188 -4584 -3178 -4583
rect -3084 -4580 -3083 -4570
rect -3081 -4580 -3080 -4570
rect -3048 -4572 -3047 -4562
rect -3045 -4572 -3044 -4562
rect -3188 -4587 -3178 -4586
rect -2968 -4647 -2967 -4627
rect -2965 -4647 -2964 -4627
rect -2925 -4681 -2924 -4670
rect -2922 -4681 -2921 -4670
rect -2968 -4702 -2967 -4682
rect -2965 -4702 -2964 -4682
rect -3137 -4827 -3136 -4807
rect -3134 -4827 -3133 -4807
rect -2609 -4798 -2604 -4792
rect -2605 -4802 -2604 -4798
rect -2602 -4796 -2601 -4792
rect -2602 -4802 -2597 -4796
rect -2790 -4836 -2789 -4826
rect -2787 -4836 -2786 -4826
rect -2854 -4846 -2853 -4836
rect -2851 -4846 -2850 -4836
rect -2821 -4846 -2820 -4836
rect -2818 -4846 -2817 -4836
rect -3094 -4861 -3093 -4850
rect -3091 -4861 -3090 -4850
rect -2609 -4852 -2604 -4846
rect -2605 -4856 -2604 -4852
rect -2602 -4850 -2601 -4846
rect -2602 -4856 -2597 -4850
rect -2587 -4850 -2586 -4846
rect -2591 -4856 -2586 -4850
rect -2584 -4850 -2583 -4846
rect -2584 -4856 -2579 -4850
rect -3137 -4882 -3136 -4862
rect -3134 -4882 -3133 -4862
rect -2937 -4914 -2932 -4908
rect -2933 -4918 -2932 -4914
rect -2930 -4912 -2929 -4908
rect -2930 -4918 -2925 -4912
rect -2937 -4968 -2932 -4962
rect -2933 -4972 -2932 -4968
rect -2930 -4966 -2929 -4962
rect -2930 -4972 -2925 -4966
rect -2915 -4966 -2914 -4962
rect -2919 -4972 -2914 -4966
rect -2912 -4966 -2911 -4962
rect -2912 -4972 -2907 -4966
<< pdiffusion >>
rect 1784 392 1785 412
rect 1787 392 1788 412
rect 1811 392 1812 412
rect 1814 392 1815 412
rect 1846 322 1847 362
rect 1849 322 1850 362
rect 2158 321 2178 322
rect 2158 318 2178 319
rect 2260 310 2261 330
rect 2263 310 2264 330
rect 2158 270 2178 271
rect 2158 267 2178 268
rect 2414 244 2415 264
rect 2417 244 2418 264
rect 2414 197 2415 216
rect 2417 197 2418 216
rect 2463 200 2464 220
rect 2466 200 2467 220
rect -3134 -2152 -3114 -2151
rect -3134 -2155 -3114 -2154
rect -3032 -2163 -3031 -2143
rect -3029 -2163 -3028 -2143
rect -3134 -2203 -3114 -2202
rect -3134 -2206 -3114 -2205
rect -2928 -2205 -2927 -2185
rect -2925 -2205 -2924 -2185
rect -2901 -2205 -2900 -2185
rect -2898 -2205 -2897 -2185
rect -2866 -2275 -2865 -2235
rect -2863 -2275 -2862 -2235
rect -2783 -2243 -2782 -2223
rect -2780 -2243 -2779 -2223
rect -2756 -2243 -2755 -2223
rect -2753 -2243 -2752 -2223
rect -2590 -2259 -2589 -2239
rect -2587 -2259 -2586 -2239
rect -2563 -2259 -2562 -2239
rect -2560 -2259 -2559 -2239
rect -2444 -2257 -2443 -2237
rect -2441 -2257 -2440 -2237
rect -2417 -2257 -2416 -2237
rect -2414 -2257 -2413 -2237
rect -2721 -2313 -2720 -2273
rect -2718 -2313 -2717 -2273
rect -2300 -2261 -2299 -2241
rect -2297 -2261 -2296 -2241
rect -2273 -2261 -2272 -2241
rect -2270 -2261 -2269 -2241
rect -2528 -2329 -2527 -2289
rect -2525 -2329 -2524 -2289
rect -2145 -2263 -2144 -2243
rect -2142 -2263 -2141 -2243
rect -2118 -2263 -2117 -2243
rect -2115 -2263 -2114 -2243
rect -3146 -2366 -3145 -2346
rect -3143 -2366 -3142 -2346
rect -3119 -2366 -3118 -2346
rect -3116 -2366 -3115 -2346
rect -2382 -2327 -2381 -2287
rect -2379 -2327 -2378 -2287
rect -2010 -2271 -2009 -2251
rect -2007 -2271 -2006 -2251
rect -1983 -2271 -1982 -2251
rect -1980 -2271 -1979 -2251
rect -2238 -2331 -2237 -2291
rect -2235 -2331 -2234 -2291
rect -2083 -2333 -2082 -2293
rect -2080 -2333 -2079 -2293
rect -1948 -2341 -1947 -2301
rect -1945 -2341 -1944 -2301
rect -1849 -2314 -1848 -2294
rect -1846 -2314 -1845 -2294
rect -1849 -2361 -1848 -2342
rect -1846 -2361 -1845 -2342
rect -3084 -2436 -3083 -2396
rect -3081 -2436 -3080 -2396
rect -1800 -2358 -1799 -2338
rect -1797 -2358 -1796 -2338
rect -1687 -2370 -1686 -2350
rect -1684 -2370 -1683 -2350
rect -1687 -2417 -1686 -2398
rect -1684 -2417 -1683 -2398
rect -1638 -2414 -1637 -2394
rect -1635 -2414 -1634 -2394
rect -1529 -2426 -1528 -2406
rect -1526 -2426 -1525 -2406
rect -1529 -2473 -1528 -2454
rect -1526 -2473 -1525 -2454
rect -1480 -2470 -1479 -2450
rect -1477 -2470 -1476 -2450
rect -1363 -2502 -1362 -2482
rect -1360 -2502 -1359 -2482
rect -1363 -2549 -1362 -2530
rect -1360 -2549 -1359 -2530
rect -1314 -2546 -1313 -2526
rect -1311 -2546 -1310 -2526
rect -3128 -3003 -3108 -3002
rect -3128 -3006 -3108 -3005
rect -3026 -3014 -3025 -2994
rect -3023 -3014 -3022 -2994
rect -2920 -3020 -2919 -3000
rect -2917 -3020 -2916 -3000
rect -2893 -3020 -2892 -3000
rect -2890 -3020 -2889 -3000
rect -2751 -3019 -2750 -2999
rect -2748 -3019 -2747 -2999
rect -2724 -3019 -2723 -2999
rect -2721 -3019 -2720 -2999
rect -2587 -3017 -2586 -2997
rect -2584 -3017 -2583 -2997
rect -2560 -3017 -2559 -2997
rect -2557 -3017 -2556 -2997
rect -2447 -3019 -2446 -2999
rect -2444 -3019 -2443 -2999
rect -2420 -3019 -2419 -2999
rect -2417 -3019 -2416 -2999
rect -2296 -3032 -2295 -3012
rect -2293 -3032 -2292 -3012
rect -2269 -3032 -2268 -3012
rect -2266 -3032 -2265 -3012
rect -3128 -3054 -3108 -3053
rect -3128 -3057 -3108 -3056
rect -2858 -3090 -2857 -3050
rect -2855 -3090 -2854 -3050
rect -2689 -3089 -2688 -3049
rect -2686 -3089 -2685 -3049
rect -2525 -3087 -2524 -3047
rect -2522 -3087 -2521 -3047
rect -2385 -3089 -2384 -3049
rect -2382 -3089 -2381 -3049
rect -1986 -3061 -1985 -3041
rect -1983 -3061 -1982 -3041
rect -2234 -3102 -2233 -3062
rect -2231 -3102 -2230 -3062
rect -1986 -3108 -1985 -3089
rect -1983 -3108 -1982 -3089
rect -1937 -3105 -1936 -3085
rect -1934 -3105 -1933 -3085
rect -2133 -3236 -2132 -3216
rect -2130 -3236 -2129 -3216
rect -2106 -3236 -2105 -3216
rect -2103 -3236 -2102 -3216
rect -3153 -3281 -3152 -3261
rect -3150 -3281 -3149 -3261
rect -3126 -3281 -3125 -3261
rect -3123 -3281 -3122 -3261
rect -2071 -3306 -2070 -3266
rect -2068 -3306 -2067 -3266
rect -1852 -3271 -1851 -3251
rect -1849 -3271 -1848 -3251
rect -3091 -3351 -3090 -3311
rect -3088 -3351 -3087 -3311
rect -1852 -3318 -1851 -3299
rect -1849 -3318 -1848 -3299
rect -1803 -3315 -1802 -3295
rect -1800 -3315 -1799 -3295
rect -1705 -3431 -1704 -3411
rect -1702 -3431 -1701 -3411
rect -1495 -3428 -1494 -3424
rect -1705 -3478 -1704 -3459
rect -1702 -3478 -1701 -3459
rect -1499 -3444 -1494 -3428
rect -1492 -3440 -1487 -3424
rect -1492 -3444 -1491 -3440
rect -1656 -3475 -1655 -3455
rect -1653 -3475 -1652 -3455
rect -1495 -3483 -1494 -3479
rect -1499 -3499 -1494 -3483
rect -1492 -3495 -1487 -3479
rect -1492 -3499 -1491 -3495
rect -1481 -3495 -1476 -3479
rect -1477 -3499 -1476 -3495
rect -1474 -3495 -1469 -3479
rect -1474 -3499 -1473 -3495
rect -3128 -3771 -3108 -3770
rect -3128 -3774 -3108 -3773
rect -3026 -3782 -3025 -3762
rect -3023 -3782 -3022 -3762
rect -2899 -3793 -2898 -3773
rect -2896 -3793 -2895 -3773
rect -2872 -3793 -2871 -3773
rect -2869 -3793 -2868 -3773
rect -3128 -3822 -3108 -3821
rect -3128 -3825 -3108 -3824
rect -2837 -3863 -2836 -3823
rect -2834 -3863 -2833 -3823
rect -2733 -3921 -2732 -3901
rect -2730 -3921 -2729 -3901
rect -2733 -3968 -2732 -3949
rect -2730 -3968 -2729 -3949
rect -2898 -3998 -2897 -3978
rect -2895 -3998 -2894 -3978
rect -2871 -3998 -2870 -3978
rect -2868 -3998 -2867 -3978
rect -2684 -3965 -2683 -3945
rect -2681 -3965 -2680 -3945
rect -2836 -4068 -2835 -4028
rect -2833 -4068 -2832 -4028
rect -2587 -4034 -2586 -4014
rect -2584 -4034 -2583 -4014
rect -2413 -4039 -2412 -4035
rect -2587 -4081 -2586 -4062
rect -2584 -4081 -2583 -4062
rect -2417 -4055 -2412 -4039
rect -2410 -4051 -2405 -4035
rect -2410 -4055 -2409 -4051
rect -2538 -4078 -2537 -4058
rect -2535 -4078 -2534 -4058
rect -2413 -4094 -2412 -4090
rect -3159 -4130 -3158 -4110
rect -3156 -4130 -3155 -4110
rect -3132 -4130 -3131 -4110
rect -3129 -4130 -3128 -4110
rect -2417 -4110 -2412 -4094
rect -2410 -4106 -2405 -4090
rect -2410 -4110 -2409 -4106
rect -2399 -4106 -2394 -4090
rect -2395 -4110 -2394 -4106
rect -2392 -4106 -2387 -4090
rect -2392 -4110 -2391 -4106
rect 712 -4139 713 -4135
rect 708 -4155 713 -4139
rect 715 -4151 720 -4135
rect 715 -4155 716 -4151
rect -3097 -4200 -3096 -4160
rect -3094 -4200 -3093 -4160
rect 712 -4194 713 -4190
rect 708 -4210 713 -4194
rect 715 -4206 720 -4190
rect 715 -4210 716 -4206
rect 726 -4206 731 -4190
rect 730 -4210 731 -4206
rect 733 -4206 738 -4190
rect 733 -4210 734 -4206
rect -3150 -4533 -3130 -4532
rect -3150 -4536 -3130 -4535
rect -3048 -4544 -3047 -4524
rect -3045 -4544 -3044 -4524
rect -2987 -4573 -2986 -4553
rect -2984 -4573 -2983 -4553
rect -2960 -4573 -2959 -4553
rect -2957 -4573 -2956 -4553
rect -3150 -4584 -3130 -4583
rect -3150 -4587 -3130 -4586
rect -2925 -4643 -2924 -4603
rect -2922 -4643 -2921 -4603
rect -3156 -4753 -3155 -4733
rect -3153 -4753 -3152 -4733
rect -3129 -4753 -3128 -4733
rect -3126 -4753 -3125 -4733
rect -2839 -4764 -2838 -4744
rect -2836 -4764 -2835 -4744
rect -2605 -4763 -2604 -4759
rect -3094 -4823 -3093 -4783
rect -3091 -4823 -3090 -4783
rect -2839 -4811 -2838 -4792
rect -2836 -4811 -2835 -4792
rect -2609 -4779 -2604 -4763
rect -2602 -4775 -2597 -4759
rect -2602 -4779 -2601 -4775
rect -2790 -4808 -2789 -4788
rect -2787 -4808 -2786 -4788
rect -2605 -4818 -2604 -4814
rect -2609 -4834 -2604 -4818
rect -2602 -4830 -2597 -4814
rect -2602 -4834 -2601 -4830
rect -2591 -4830 -2586 -4814
rect -2587 -4834 -2586 -4830
rect -2584 -4830 -2579 -4814
rect -2584 -4834 -2583 -4830
rect -2933 -4879 -2932 -4875
rect -2937 -4895 -2932 -4879
rect -2930 -4891 -2925 -4875
rect -2930 -4895 -2929 -4891
rect -2933 -4934 -2932 -4930
rect -2937 -4950 -2932 -4934
rect -2930 -4946 -2925 -4930
rect -2930 -4950 -2929 -4946
rect -2919 -4946 -2914 -4930
rect -2915 -4950 -2914 -4946
rect -2912 -4946 -2907 -4930
rect -2912 -4950 -2911 -4946
<< ndcontact >>
rect 1799 318 1803 338
rect 1807 318 1811 338
rect 2120 322 2130 326
rect 2120 314 2130 318
rect 2220 307 2224 317
rect 2228 307 2232 317
rect 1842 284 1846 295
rect 1850 284 1854 295
rect 1799 263 1803 283
rect 1807 263 1811 283
rect 2120 271 2130 275
rect 2220 274 2224 284
rect 2228 274 2232 284
rect 2256 282 2260 292
rect 2264 282 2268 292
rect 2120 263 2130 267
rect 2459 172 2463 182
rect 2467 172 2471 182
rect 2395 162 2399 172
rect 2403 162 2407 172
rect 2428 162 2432 172
rect 2436 162 2440 172
rect -3172 -2151 -3162 -2147
rect -3172 -2159 -3162 -2155
rect -3072 -2166 -3068 -2158
rect -3064 -2166 -3060 -2158
rect -3172 -2202 -3162 -2198
rect -3072 -2199 -3068 -2189
rect -3064 -2199 -3060 -2189
rect -3036 -2191 -3032 -2181
rect -3028 -2191 -3024 -2181
rect -3172 -2210 -3162 -2206
rect -2913 -2279 -2909 -2259
rect -2905 -2279 -2901 -2259
rect -2870 -2313 -2866 -2302
rect -2862 -2313 -2858 -2302
rect -2913 -2334 -2909 -2314
rect -2905 -2334 -2901 -2314
rect -2768 -2317 -2764 -2297
rect -2760 -2317 -2756 -2297
rect -2575 -2333 -2571 -2313
rect -2567 -2333 -2563 -2313
rect -2725 -2351 -2721 -2340
rect -2717 -2351 -2713 -2340
rect -2768 -2372 -2764 -2352
rect -2760 -2372 -2756 -2352
rect -2429 -2331 -2425 -2311
rect -2421 -2331 -2417 -2311
rect -2285 -2335 -2281 -2315
rect -2277 -2335 -2273 -2315
rect -2532 -2367 -2528 -2356
rect -2524 -2367 -2520 -2356
rect -2386 -2365 -2382 -2354
rect -2378 -2365 -2374 -2354
rect -2130 -2337 -2126 -2317
rect -2122 -2337 -2118 -2317
rect -2575 -2388 -2571 -2368
rect -2567 -2388 -2563 -2368
rect -2429 -2386 -2425 -2366
rect -2421 -2386 -2417 -2366
rect -2242 -2369 -2238 -2358
rect -2234 -2369 -2230 -2358
rect -1995 -2345 -1991 -2325
rect -1987 -2345 -1983 -2325
rect -2285 -2390 -2281 -2370
rect -2277 -2390 -2273 -2370
rect -2087 -2371 -2083 -2360
rect -2079 -2371 -2075 -2360
rect -2130 -2392 -2126 -2372
rect -2122 -2392 -2118 -2372
rect -1952 -2379 -1948 -2368
rect -1944 -2379 -1940 -2368
rect -3131 -2440 -3127 -2420
rect -3123 -2440 -3119 -2420
rect -1995 -2400 -1991 -2380
rect -1987 -2400 -1983 -2380
rect -1804 -2386 -1800 -2376
rect -1796 -2386 -1792 -2376
rect -1868 -2396 -1864 -2386
rect -1860 -2396 -1856 -2386
rect -1835 -2396 -1831 -2386
rect -1827 -2396 -1823 -2386
rect -1642 -2442 -1638 -2432
rect -1634 -2442 -1630 -2432
rect -1706 -2452 -1702 -2442
rect -1698 -2452 -1694 -2442
rect -1673 -2452 -1669 -2442
rect -1665 -2452 -1661 -2442
rect -3088 -2474 -3084 -2463
rect -3080 -2474 -3076 -2463
rect -3131 -2495 -3127 -2475
rect -3123 -2495 -3119 -2475
rect -1484 -2498 -1480 -2488
rect -1476 -2498 -1472 -2488
rect -1548 -2508 -1544 -2498
rect -1540 -2508 -1536 -2498
rect -1515 -2508 -1511 -2498
rect -1507 -2508 -1503 -2498
rect -1318 -2574 -1314 -2564
rect -1310 -2574 -1306 -2564
rect -1382 -2584 -1378 -2574
rect -1374 -2584 -1370 -2574
rect -1349 -2584 -1345 -2574
rect -1341 -2584 -1337 -2574
rect -3166 -3002 -3156 -2998
rect -3166 -3010 -3156 -3006
rect -3066 -3017 -3062 -3009
rect -3058 -3017 -3054 -3009
rect -3166 -3053 -3156 -3049
rect -3066 -3050 -3062 -3040
rect -3058 -3050 -3054 -3040
rect -3030 -3042 -3026 -3032
rect -3022 -3042 -3018 -3032
rect -3166 -3061 -3156 -3057
rect -2905 -3094 -2901 -3074
rect -2897 -3094 -2893 -3074
rect -2736 -3093 -2732 -3073
rect -2728 -3093 -2724 -3073
rect -2572 -3091 -2568 -3071
rect -2564 -3091 -2560 -3071
rect -2432 -3093 -2428 -3073
rect -2424 -3093 -2420 -3073
rect -2862 -3128 -2858 -3117
rect -2854 -3128 -2850 -3117
rect -2693 -3127 -2689 -3116
rect -2685 -3127 -2681 -3116
rect -2529 -3125 -2525 -3114
rect -2521 -3125 -2517 -3114
rect -2281 -3106 -2277 -3086
rect -2273 -3106 -2269 -3086
rect -2905 -3149 -2901 -3129
rect -2897 -3149 -2893 -3129
rect -2736 -3148 -2732 -3128
rect -2728 -3148 -2724 -3128
rect -2572 -3146 -2568 -3126
rect -2564 -3146 -2560 -3126
rect -2389 -3127 -2385 -3116
rect -2381 -3127 -2377 -3116
rect -2432 -3148 -2428 -3128
rect -2424 -3148 -2420 -3128
rect -2238 -3140 -2234 -3129
rect -2230 -3140 -2226 -3129
rect -1941 -3133 -1937 -3123
rect -1933 -3133 -1929 -3123
rect -2281 -3161 -2277 -3141
rect -2273 -3161 -2269 -3141
rect -2005 -3143 -2001 -3133
rect -1997 -3143 -1993 -3133
rect -1972 -3143 -1968 -3133
rect -1964 -3143 -1960 -3133
rect -2118 -3310 -2114 -3290
rect -2110 -3310 -2106 -3290
rect -3138 -3355 -3134 -3335
rect -3130 -3355 -3126 -3335
rect -2075 -3344 -2071 -3333
rect -2067 -3344 -2063 -3333
rect -1807 -3343 -1803 -3333
rect -1799 -3343 -1795 -3333
rect -2118 -3365 -2114 -3345
rect -2110 -3365 -2106 -3345
rect -1871 -3353 -1867 -3343
rect -1863 -3353 -1859 -3343
rect -1838 -3353 -1834 -3343
rect -1830 -3353 -1826 -3343
rect -3095 -3389 -3091 -3378
rect -3087 -3389 -3083 -3378
rect -3138 -3410 -3134 -3390
rect -3130 -3410 -3126 -3390
rect -1499 -3467 -1495 -3463
rect -1491 -3461 -1487 -3457
rect -1660 -3503 -1656 -3493
rect -1652 -3503 -1648 -3493
rect -1724 -3513 -1720 -3503
rect -1716 -3513 -1712 -3503
rect -1691 -3513 -1687 -3503
rect -1683 -3513 -1679 -3503
rect -1499 -3521 -1495 -3517
rect -1491 -3515 -1487 -3511
rect -1481 -3515 -1477 -3511
rect -1473 -3515 -1469 -3511
rect -3166 -3770 -3156 -3766
rect -3166 -3778 -3156 -3774
rect -3066 -3785 -3062 -3777
rect -3058 -3785 -3054 -3777
rect -3166 -3821 -3156 -3817
rect -3066 -3818 -3062 -3808
rect -3058 -3818 -3054 -3808
rect -3030 -3810 -3026 -3800
rect -3022 -3810 -3018 -3800
rect -3166 -3829 -3156 -3825
rect -2884 -3867 -2880 -3847
rect -2876 -3867 -2872 -3847
rect -2841 -3901 -2837 -3890
rect -2833 -3901 -2829 -3890
rect -2884 -3922 -2880 -3902
rect -2876 -3922 -2872 -3902
rect -2688 -3993 -2684 -3983
rect -2680 -3993 -2676 -3983
rect -2752 -4003 -2748 -3993
rect -2744 -4003 -2740 -3993
rect -2719 -4003 -2715 -3993
rect -2711 -4003 -2707 -3993
rect -2883 -4072 -2879 -4052
rect -2875 -4072 -2871 -4052
rect -2840 -4106 -2836 -4095
rect -2832 -4106 -2828 -4095
rect -2417 -4078 -2413 -4074
rect -2409 -4072 -2405 -4068
rect -2542 -4106 -2538 -4096
rect -2534 -4106 -2530 -4096
rect -2883 -4127 -2879 -4107
rect -2875 -4127 -2871 -4107
rect -2606 -4116 -2602 -4106
rect -2598 -4116 -2594 -4106
rect -2573 -4116 -2569 -4106
rect -2565 -4116 -2561 -4106
rect -2417 -4132 -2413 -4128
rect -2409 -4126 -2405 -4122
rect -2399 -4126 -2395 -4122
rect -2391 -4126 -2387 -4122
rect -3144 -4204 -3140 -4184
rect -3136 -4204 -3132 -4184
rect 708 -4178 712 -4174
rect 716 -4172 720 -4168
rect -3101 -4238 -3097 -4227
rect -3093 -4238 -3089 -4227
rect 708 -4232 712 -4228
rect 716 -4226 720 -4222
rect 726 -4226 730 -4222
rect 734 -4226 738 -4222
rect -3144 -4259 -3140 -4239
rect -3136 -4259 -3132 -4239
rect -3188 -4532 -3178 -4528
rect -3188 -4540 -3178 -4536
rect -3088 -4547 -3084 -4539
rect -3080 -4547 -3076 -4539
rect -3188 -4583 -3178 -4579
rect -3088 -4580 -3084 -4570
rect -3080 -4580 -3076 -4570
rect -3052 -4572 -3048 -4562
rect -3044 -4572 -3040 -4562
rect -3188 -4591 -3178 -4587
rect -2972 -4647 -2968 -4627
rect -2964 -4647 -2960 -4627
rect -2929 -4681 -2925 -4670
rect -2921 -4681 -2917 -4670
rect -2972 -4702 -2968 -4682
rect -2964 -4702 -2960 -4682
rect -3141 -4827 -3137 -4807
rect -3133 -4827 -3129 -4807
rect -2609 -4802 -2605 -4798
rect -2601 -4796 -2597 -4792
rect -2794 -4836 -2790 -4826
rect -2786 -4836 -2782 -4826
rect -2858 -4846 -2854 -4836
rect -2850 -4846 -2846 -4836
rect -2825 -4846 -2821 -4836
rect -2817 -4846 -2813 -4836
rect -3098 -4861 -3094 -4850
rect -3090 -4861 -3086 -4850
rect -2609 -4856 -2605 -4852
rect -2601 -4850 -2597 -4846
rect -2591 -4850 -2587 -4846
rect -2583 -4850 -2579 -4846
rect -3141 -4882 -3137 -4862
rect -3133 -4882 -3129 -4862
rect -2937 -4918 -2933 -4914
rect -2929 -4912 -2925 -4908
rect -2937 -4972 -2933 -4968
rect -2929 -4966 -2925 -4962
rect -2919 -4966 -2915 -4962
rect -2911 -4966 -2907 -4962
<< pdcontact >>
rect 1780 392 1784 412
rect 1788 392 1792 412
rect 1807 392 1811 412
rect 1815 392 1819 412
rect 1842 322 1846 362
rect 1850 322 1854 362
rect 2158 322 2178 326
rect 2158 314 2178 318
rect 2256 310 2260 330
rect 2264 310 2268 330
rect 2158 271 2178 275
rect 2158 263 2178 267
rect 2410 244 2414 264
rect 2418 244 2422 264
rect 2410 197 2414 216
rect 2418 197 2422 216
rect 2459 200 2463 220
rect 2467 200 2471 220
rect -3134 -2151 -3114 -2147
rect -3134 -2159 -3114 -2155
rect -3036 -2163 -3032 -2143
rect -3028 -2163 -3024 -2143
rect -3134 -2202 -3114 -2198
rect -2932 -2205 -2928 -2185
rect -2924 -2205 -2920 -2185
rect -2905 -2205 -2901 -2185
rect -2897 -2205 -2893 -2185
rect -3134 -2210 -3114 -2206
rect -2870 -2275 -2866 -2235
rect -2862 -2275 -2858 -2235
rect -2787 -2243 -2783 -2223
rect -2779 -2243 -2775 -2223
rect -2760 -2243 -2756 -2223
rect -2752 -2243 -2748 -2223
rect -2594 -2259 -2590 -2239
rect -2586 -2259 -2582 -2239
rect -2567 -2259 -2563 -2239
rect -2559 -2259 -2555 -2239
rect -2448 -2257 -2444 -2237
rect -2440 -2257 -2436 -2237
rect -2421 -2257 -2417 -2237
rect -2413 -2257 -2409 -2237
rect -2725 -2313 -2721 -2273
rect -2717 -2313 -2713 -2273
rect -2304 -2261 -2300 -2241
rect -2296 -2261 -2292 -2241
rect -2277 -2261 -2273 -2241
rect -2269 -2261 -2265 -2241
rect -2532 -2329 -2528 -2289
rect -2524 -2329 -2520 -2289
rect -2149 -2263 -2145 -2243
rect -2141 -2263 -2137 -2243
rect -2122 -2263 -2118 -2243
rect -2114 -2263 -2110 -2243
rect -3150 -2366 -3146 -2346
rect -3142 -2366 -3138 -2346
rect -3123 -2366 -3119 -2346
rect -3115 -2366 -3111 -2346
rect -2386 -2327 -2382 -2287
rect -2378 -2327 -2374 -2287
rect -2014 -2271 -2010 -2251
rect -2006 -2271 -2002 -2251
rect -1987 -2271 -1983 -2251
rect -1979 -2271 -1975 -2251
rect -2242 -2331 -2238 -2291
rect -2234 -2331 -2230 -2291
rect -2087 -2333 -2083 -2293
rect -2079 -2333 -2075 -2293
rect -1952 -2341 -1948 -2301
rect -1944 -2341 -1940 -2301
rect -1853 -2314 -1849 -2294
rect -1845 -2314 -1841 -2294
rect -1853 -2361 -1849 -2342
rect -1845 -2361 -1841 -2342
rect -3088 -2436 -3084 -2396
rect -3080 -2436 -3076 -2396
rect -1804 -2358 -1800 -2338
rect -1796 -2358 -1792 -2338
rect -1691 -2370 -1687 -2350
rect -1683 -2370 -1679 -2350
rect -1691 -2417 -1687 -2398
rect -1683 -2417 -1679 -2398
rect -1642 -2414 -1638 -2394
rect -1634 -2414 -1630 -2394
rect -1533 -2426 -1529 -2406
rect -1525 -2426 -1521 -2406
rect -1533 -2473 -1529 -2454
rect -1525 -2473 -1521 -2454
rect -1484 -2470 -1480 -2450
rect -1476 -2470 -1472 -2450
rect -1367 -2502 -1363 -2482
rect -1359 -2502 -1355 -2482
rect -1367 -2549 -1363 -2530
rect -1359 -2549 -1355 -2530
rect -1318 -2546 -1314 -2526
rect -1310 -2546 -1306 -2526
rect -3128 -3002 -3108 -2998
rect -3128 -3010 -3108 -3006
rect -3030 -3014 -3026 -2994
rect -3022 -3014 -3018 -2994
rect -2924 -3020 -2920 -3000
rect -2916 -3020 -2912 -3000
rect -2897 -3020 -2893 -3000
rect -2889 -3020 -2885 -3000
rect -2755 -3019 -2751 -2999
rect -2747 -3019 -2743 -2999
rect -2728 -3019 -2724 -2999
rect -2720 -3019 -2716 -2999
rect -2591 -3017 -2587 -2997
rect -2583 -3017 -2579 -2997
rect -2564 -3017 -2560 -2997
rect -2556 -3017 -2552 -2997
rect -3128 -3053 -3108 -3049
rect -2451 -3019 -2447 -2999
rect -2443 -3019 -2439 -2999
rect -2424 -3019 -2420 -2999
rect -2416 -3019 -2412 -2999
rect -2300 -3032 -2296 -3012
rect -2292 -3032 -2288 -3012
rect -2273 -3032 -2269 -3012
rect -2265 -3032 -2261 -3012
rect -3128 -3061 -3108 -3057
rect -2862 -3090 -2858 -3050
rect -2854 -3090 -2850 -3050
rect -2693 -3089 -2689 -3049
rect -2685 -3089 -2681 -3049
rect -2529 -3087 -2525 -3047
rect -2521 -3087 -2517 -3047
rect -2389 -3089 -2385 -3049
rect -2381 -3089 -2377 -3049
rect -1990 -3061 -1986 -3041
rect -1982 -3061 -1978 -3041
rect -2238 -3102 -2234 -3062
rect -2230 -3102 -2226 -3062
rect -1990 -3108 -1986 -3089
rect -1982 -3108 -1978 -3089
rect -1941 -3105 -1937 -3085
rect -1933 -3105 -1929 -3085
rect -2137 -3236 -2133 -3216
rect -2129 -3236 -2125 -3216
rect -2110 -3236 -2106 -3216
rect -2102 -3236 -2098 -3216
rect -3157 -3281 -3153 -3261
rect -3149 -3281 -3145 -3261
rect -3130 -3281 -3126 -3261
rect -3122 -3281 -3118 -3261
rect -2075 -3306 -2071 -3266
rect -2067 -3306 -2063 -3266
rect -1856 -3271 -1852 -3251
rect -1848 -3271 -1844 -3251
rect -3095 -3351 -3091 -3311
rect -3087 -3351 -3083 -3311
rect -1856 -3318 -1852 -3299
rect -1848 -3318 -1844 -3299
rect -1807 -3315 -1803 -3295
rect -1799 -3315 -1795 -3295
rect -1709 -3431 -1705 -3411
rect -1701 -3431 -1697 -3411
rect -1499 -3428 -1495 -3424
rect -1709 -3478 -1705 -3459
rect -1701 -3478 -1697 -3459
rect -1491 -3444 -1487 -3440
rect -1660 -3475 -1656 -3455
rect -1652 -3475 -1648 -3455
rect -1499 -3483 -1495 -3479
rect -1491 -3499 -1487 -3495
rect -1481 -3499 -1477 -3495
rect -1473 -3499 -1469 -3495
rect -3128 -3770 -3108 -3766
rect -3128 -3778 -3108 -3774
rect -3030 -3782 -3026 -3762
rect -3022 -3782 -3018 -3762
rect -2903 -3793 -2899 -3773
rect -2895 -3793 -2891 -3773
rect -2876 -3793 -2872 -3773
rect -2868 -3793 -2864 -3773
rect -3128 -3821 -3108 -3817
rect -3128 -3829 -3108 -3825
rect -2841 -3863 -2837 -3823
rect -2833 -3863 -2829 -3823
rect -2737 -3921 -2733 -3901
rect -2729 -3921 -2725 -3901
rect -2737 -3968 -2733 -3949
rect -2729 -3968 -2725 -3949
rect -2902 -3998 -2898 -3978
rect -2894 -3998 -2890 -3978
rect -2875 -3998 -2871 -3978
rect -2867 -3998 -2863 -3978
rect -2688 -3965 -2684 -3945
rect -2680 -3965 -2676 -3945
rect -2840 -4068 -2836 -4028
rect -2832 -4068 -2828 -4028
rect -2591 -4034 -2587 -4014
rect -2583 -4034 -2579 -4014
rect -2417 -4039 -2413 -4035
rect -2591 -4081 -2587 -4062
rect -2583 -4081 -2579 -4062
rect -2409 -4055 -2405 -4051
rect -2542 -4078 -2538 -4058
rect -2534 -4078 -2530 -4058
rect -2417 -4094 -2413 -4090
rect -3163 -4130 -3159 -4110
rect -3155 -4130 -3151 -4110
rect -3136 -4130 -3132 -4110
rect -3128 -4130 -3124 -4110
rect -2409 -4110 -2405 -4106
rect -2399 -4110 -2395 -4106
rect -2391 -4110 -2387 -4106
rect 708 -4139 712 -4135
rect 716 -4155 720 -4151
rect -3101 -4200 -3097 -4160
rect -3093 -4200 -3089 -4160
rect 708 -4194 712 -4190
rect 716 -4210 720 -4206
rect 726 -4210 730 -4206
rect 734 -4210 738 -4206
rect -3150 -4532 -3130 -4528
rect -3150 -4540 -3130 -4536
rect -3052 -4544 -3048 -4524
rect -3044 -4544 -3040 -4524
rect -3150 -4583 -3130 -4579
rect -2991 -4573 -2987 -4553
rect -2983 -4573 -2979 -4553
rect -2964 -4573 -2960 -4553
rect -2956 -4573 -2952 -4553
rect -3150 -4591 -3130 -4587
rect -2929 -4643 -2925 -4603
rect -2921 -4643 -2917 -4603
rect -3160 -4753 -3156 -4733
rect -3152 -4753 -3148 -4733
rect -3133 -4753 -3129 -4733
rect -3125 -4753 -3121 -4733
rect -2843 -4764 -2839 -4744
rect -2835 -4764 -2831 -4744
rect -2609 -4763 -2605 -4759
rect -3098 -4823 -3094 -4783
rect -3090 -4823 -3086 -4783
rect -2843 -4811 -2839 -4792
rect -2835 -4811 -2831 -4792
rect -2601 -4779 -2597 -4775
rect -2794 -4808 -2790 -4788
rect -2786 -4808 -2782 -4788
rect -2609 -4818 -2605 -4814
rect -2601 -4834 -2597 -4830
rect -2591 -4834 -2587 -4830
rect -2583 -4834 -2579 -4830
rect -2937 -4879 -2933 -4875
rect -2929 -4895 -2925 -4891
rect -2937 -4934 -2933 -4930
rect -2929 -4950 -2925 -4946
rect -2919 -4950 -2915 -4946
rect -2911 -4950 -2907 -4946
<< psubstratepcontact >>
rect 2109 329 2113 333
rect 2109 308 2113 312
rect 2109 278 2113 282
rect 1835 273 1839 277
rect 1856 273 1860 277
rect 2249 267 2253 271
rect 2270 267 2274 271
rect 2109 257 2113 261
rect 1792 252 1796 256
rect 1813 252 1817 256
rect 2452 157 2456 161
rect 2473 157 2477 161
rect 2388 150 2392 154
rect 2409 150 2413 154
rect 2421 150 2425 154
rect 2442 150 2446 154
rect -3183 -2144 -3179 -2140
rect -3183 -2165 -3179 -2161
rect -3183 -2195 -3179 -2191
rect -3043 -2206 -3039 -2202
rect -3022 -2206 -3018 -2202
rect -3183 -2216 -3179 -2212
rect -2877 -2324 -2873 -2320
rect -2856 -2324 -2852 -2320
rect -2920 -2345 -2916 -2341
rect -2899 -2345 -2895 -2341
rect -2732 -2362 -2728 -2358
rect -2711 -2362 -2707 -2358
rect -2775 -2383 -2771 -2379
rect -2754 -2383 -2750 -2379
rect -2539 -2378 -2535 -2374
rect -2518 -2378 -2514 -2374
rect -2393 -2376 -2389 -2372
rect -2372 -2376 -2368 -2372
rect -2249 -2380 -2245 -2376
rect -2228 -2380 -2224 -2376
rect -2094 -2382 -2090 -2378
rect -2073 -2382 -2069 -2378
rect -2582 -2399 -2578 -2395
rect -2561 -2399 -2557 -2395
rect -2436 -2397 -2432 -2393
rect -2415 -2397 -2411 -2393
rect -2292 -2401 -2288 -2397
rect -2271 -2401 -2267 -2397
rect -2137 -2403 -2133 -2399
rect -2116 -2403 -2112 -2399
rect -1959 -2390 -1955 -2386
rect -1938 -2390 -1934 -2386
rect -1811 -2401 -1807 -2397
rect -1790 -2401 -1786 -2397
rect -2002 -2411 -1998 -2407
rect -1981 -2411 -1977 -2407
rect -1875 -2408 -1871 -2404
rect -1854 -2408 -1850 -2404
rect -1842 -2408 -1838 -2404
rect -1821 -2408 -1817 -2404
rect -1649 -2457 -1645 -2453
rect -1628 -2457 -1624 -2453
rect -1713 -2464 -1709 -2460
rect -1692 -2464 -1688 -2460
rect -1680 -2464 -1676 -2460
rect -1659 -2464 -1655 -2460
rect -3095 -2485 -3091 -2481
rect -3074 -2485 -3070 -2481
rect -3138 -2506 -3134 -2502
rect -3117 -2506 -3113 -2502
rect -1491 -2513 -1487 -2509
rect -1470 -2513 -1466 -2509
rect -1555 -2520 -1551 -2516
rect -1534 -2520 -1530 -2516
rect -1522 -2520 -1518 -2516
rect -1501 -2520 -1497 -2516
rect -1325 -2589 -1321 -2585
rect -1304 -2589 -1300 -2585
rect -1389 -2596 -1385 -2592
rect -1368 -2596 -1364 -2592
rect -1356 -2596 -1352 -2592
rect -1335 -2596 -1331 -2592
rect -3177 -2995 -3173 -2991
rect -3177 -3016 -3173 -3012
rect -3177 -3046 -3173 -3042
rect -3037 -3057 -3033 -3053
rect -3016 -3057 -3012 -3053
rect -3177 -3067 -3173 -3063
rect -2869 -3139 -2865 -3135
rect -2848 -3139 -2844 -3135
rect -2700 -3138 -2696 -3134
rect -2679 -3138 -2675 -3134
rect -2536 -3136 -2532 -3132
rect -2515 -3136 -2511 -3132
rect -2396 -3138 -2392 -3134
rect -2375 -3138 -2371 -3134
rect -2912 -3160 -2908 -3156
rect -2891 -3160 -2887 -3156
rect -2743 -3159 -2739 -3155
rect -2722 -3159 -2718 -3155
rect -2579 -3157 -2575 -3153
rect -2558 -3157 -2554 -3153
rect -2439 -3159 -2435 -3155
rect -2418 -3159 -2414 -3155
rect -2245 -3151 -2241 -3147
rect -2224 -3151 -2220 -3147
rect -1948 -3148 -1944 -3144
rect -1927 -3148 -1923 -3144
rect -2012 -3155 -2008 -3151
rect -1991 -3155 -1987 -3151
rect -1979 -3155 -1975 -3151
rect -1958 -3155 -1954 -3151
rect -2288 -3172 -2284 -3168
rect -2267 -3172 -2263 -3168
rect -2082 -3355 -2078 -3351
rect -2061 -3355 -2057 -3351
rect -1814 -3358 -1810 -3354
rect -1793 -3358 -1789 -3354
rect -1878 -3365 -1874 -3361
rect -1857 -3365 -1853 -3361
rect -1845 -3365 -1841 -3361
rect -1824 -3365 -1820 -3361
rect -2125 -3376 -2121 -3372
rect -2104 -3376 -2100 -3372
rect -3102 -3400 -3098 -3396
rect -3081 -3400 -3077 -3396
rect -3145 -3421 -3141 -3417
rect -3124 -3421 -3120 -3417
rect -1667 -3518 -1663 -3514
rect -1646 -3518 -1642 -3514
rect -1731 -3525 -1727 -3521
rect -1710 -3525 -1706 -3521
rect -1698 -3525 -1694 -3521
rect -1677 -3525 -1673 -3521
rect -3177 -3763 -3173 -3759
rect -3177 -3784 -3173 -3780
rect -3177 -3814 -3173 -3810
rect -3037 -3825 -3033 -3821
rect -3016 -3825 -3012 -3821
rect -3177 -3835 -3173 -3831
rect -2848 -3912 -2844 -3908
rect -2827 -3912 -2823 -3908
rect -2891 -3933 -2887 -3929
rect -2870 -3933 -2866 -3929
rect -2695 -4008 -2691 -4004
rect -2674 -4008 -2670 -4004
rect -2759 -4015 -2755 -4011
rect -2738 -4015 -2734 -4011
rect -2726 -4015 -2722 -4011
rect -2705 -4015 -2701 -4011
rect -2847 -4117 -2843 -4113
rect -2826 -4117 -2822 -4113
rect -2549 -4121 -2545 -4117
rect -2528 -4121 -2524 -4117
rect -2613 -4128 -2609 -4124
rect -2592 -4128 -2588 -4124
rect -2580 -4128 -2576 -4124
rect -2559 -4128 -2555 -4124
rect -2890 -4138 -2886 -4134
rect -2869 -4138 -2865 -4134
rect -3108 -4249 -3104 -4245
rect -3087 -4249 -3083 -4245
rect -3151 -4270 -3147 -4266
rect -3130 -4270 -3126 -4266
rect -3199 -4525 -3195 -4521
rect -3199 -4546 -3195 -4542
rect -3199 -4576 -3195 -4572
rect -3059 -4587 -3055 -4583
rect -3038 -4587 -3034 -4583
rect -3199 -4597 -3195 -4593
rect -2936 -4692 -2932 -4688
rect -2915 -4692 -2911 -4688
rect -2979 -4713 -2975 -4709
rect -2958 -4713 -2954 -4709
rect -2801 -4851 -2797 -4847
rect -2780 -4851 -2776 -4847
rect -2865 -4858 -2861 -4854
rect -2844 -4858 -2840 -4854
rect -2832 -4858 -2828 -4854
rect -2811 -4858 -2807 -4854
rect -3105 -4872 -3101 -4868
rect -3084 -4872 -3080 -4868
rect -3148 -4893 -3144 -4889
rect -3127 -4893 -3123 -4889
<< nsubstratencontact >>
rect 1775 439 1779 443
rect 1792 439 1796 443
rect 1802 439 1806 443
rect 1819 439 1823 443
rect 1837 369 1841 373
rect 1854 369 1858 373
rect 2195 327 2199 331
rect 2251 340 2255 344
rect 2268 340 2272 344
rect 2195 310 2199 314
rect 2195 276 2199 280
rect 2405 278 2409 282
rect 2422 278 2426 282
rect 2195 259 2199 263
rect 2454 230 2458 234
rect 2471 230 2475 234
rect -3097 -2146 -3093 -2142
rect -3041 -2133 -3037 -2129
rect -3024 -2133 -3020 -2129
rect -3097 -2163 -3093 -2159
rect -2937 -2158 -2933 -2154
rect -2920 -2158 -2916 -2154
rect -2910 -2158 -2906 -2154
rect -2893 -2158 -2889 -2154
rect -3097 -2197 -3093 -2193
rect -2792 -2196 -2788 -2192
rect -2775 -2196 -2771 -2192
rect -2765 -2196 -2761 -2192
rect -2748 -2196 -2744 -2192
rect -3097 -2214 -3093 -2210
rect -2599 -2212 -2595 -2208
rect -2582 -2212 -2578 -2208
rect -2572 -2212 -2568 -2208
rect -2555 -2212 -2551 -2208
rect -2453 -2210 -2449 -2206
rect -2436 -2210 -2432 -2206
rect -2426 -2210 -2422 -2206
rect -2409 -2210 -2405 -2206
rect -2309 -2214 -2305 -2210
rect -2292 -2214 -2288 -2210
rect -2282 -2214 -2278 -2210
rect -2265 -2214 -2261 -2210
rect -2154 -2216 -2150 -2212
rect -2137 -2216 -2133 -2212
rect -2127 -2216 -2123 -2212
rect -2110 -2216 -2106 -2212
rect -2875 -2228 -2871 -2224
rect -2858 -2228 -2854 -2224
rect -2019 -2224 -2015 -2220
rect -2002 -2224 -1998 -2220
rect -1992 -2224 -1988 -2220
rect -1975 -2224 -1971 -2220
rect -2730 -2266 -2726 -2262
rect -2713 -2266 -2709 -2262
rect -3155 -2319 -3151 -2315
rect -3138 -2319 -3134 -2315
rect -3128 -2319 -3124 -2315
rect -3111 -2319 -3107 -2315
rect -2537 -2282 -2533 -2278
rect -2520 -2282 -2516 -2278
rect -2391 -2280 -2387 -2276
rect -2374 -2280 -2370 -2276
rect -2247 -2284 -2243 -2280
rect -2230 -2284 -2226 -2280
rect -2092 -2286 -2088 -2282
rect -2075 -2286 -2071 -2282
rect -1858 -2280 -1854 -2276
rect -1841 -2280 -1837 -2276
rect -1957 -2294 -1953 -2290
rect -1940 -2294 -1936 -2290
rect -3093 -2389 -3089 -2385
rect -3076 -2389 -3072 -2385
rect -1809 -2328 -1805 -2324
rect -1792 -2328 -1788 -2324
rect -1696 -2336 -1692 -2332
rect -1679 -2336 -1675 -2332
rect -1647 -2384 -1643 -2380
rect -1630 -2384 -1626 -2380
rect -1538 -2392 -1534 -2388
rect -1521 -2392 -1517 -2388
rect -1489 -2440 -1485 -2436
rect -1472 -2440 -1468 -2436
rect -1372 -2468 -1368 -2464
rect -1355 -2468 -1351 -2464
rect -1323 -2516 -1319 -2512
rect -1306 -2516 -1302 -2512
rect -2929 -2973 -2925 -2969
rect -2912 -2973 -2908 -2969
rect -2902 -2973 -2898 -2969
rect -2885 -2973 -2881 -2969
rect -2760 -2972 -2756 -2968
rect -2743 -2972 -2739 -2968
rect -2733 -2972 -2729 -2968
rect -2716 -2972 -2712 -2968
rect -2596 -2970 -2592 -2966
rect -2579 -2970 -2575 -2966
rect -2569 -2970 -2565 -2966
rect -2552 -2970 -2548 -2966
rect -2456 -2972 -2452 -2968
rect -2439 -2972 -2435 -2968
rect -2429 -2972 -2425 -2968
rect -2412 -2972 -2408 -2968
rect -3091 -2997 -3087 -2993
rect -3035 -2984 -3031 -2980
rect -3018 -2984 -3014 -2980
rect -2305 -2985 -2301 -2981
rect -2288 -2985 -2284 -2981
rect -2278 -2985 -2274 -2981
rect -2261 -2985 -2257 -2981
rect -3091 -3014 -3087 -3010
rect -3091 -3048 -3087 -3044
rect -2867 -3043 -2863 -3039
rect -2850 -3043 -2846 -3039
rect -2698 -3042 -2694 -3038
rect -2681 -3042 -2677 -3038
rect -2534 -3040 -2530 -3036
rect -2517 -3040 -2513 -3036
rect -1995 -3027 -1991 -3023
rect -1978 -3027 -1974 -3023
rect -2394 -3042 -2390 -3038
rect -2377 -3042 -2373 -3038
rect -3091 -3065 -3087 -3061
rect -2243 -3055 -2239 -3051
rect -2226 -3055 -2222 -3051
rect -1946 -3075 -1942 -3071
rect -1929 -3075 -1925 -3071
rect -2142 -3189 -2138 -3185
rect -2125 -3189 -2121 -3185
rect -2115 -3189 -2111 -3185
rect -2098 -3189 -2094 -3185
rect -3162 -3234 -3158 -3230
rect -3145 -3234 -3141 -3230
rect -3135 -3234 -3131 -3230
rect -3118 -3234 -3114 -3230
rect -1861 -3237 -1857 -3233
rect -1844 -3237 -1840 -3233
rect -2080 -3259 -2076 -3255
rect -2063 -3259 -2059 -3255
rect -3100 -3304 -3096 -3300
rect -3083 -3304 -3079 -3300
rect -1812 -3285 -1808 -3281
rect -1795 -3285 -1791 -3281
rect -1714 -3397 -1710 -3393
rect -1697 -3397 -1693 -3393
rect -1665 -3445 -1661 -3441
rect -1648 -3445 -1644 -3441
rect -2908 -3746 -2904 -3742
rect -2891 -3746 -2887 -3742
rect -2881 -3746 -2877 -3742
rect -2864 -3746 -2860 -3742
rect -3091 -3765 -3087 -3761
rect -3035 -3752 -3031 -3748
rect -3018 -3752 -3014 -3748
rect -3091 -3782 -3087 -3778
rect -3091 -3816 -3087 -3812
rect -2846 -3816 -2842 -3812
rect -2829 -3816 -2825 -3812
rect -3091 -3833 -3087 -3829
rect -2742 -3887 -2738 -3883
rect -2725 -3887 -2721 -3883
rect -2907 -3951 -2903 -3947
rect -2890 -3951 -2886 -3947
rect -2880 -3951 -2876 -3947
rect -2863 -3951 -2859 -3947
rect -2693 -3935 -2689 -3931
rect -2676 -3935 -2672 -3931
rect -2596 -4000 -2592 -3996
rect -2579 -4000 -2575 -3996
rect -2845 -4021 -2841 -4017
rect -2828 -4021 -2824 -4017
rect -3168 -4083 -3164 -4079
rect -3151 -4083 -3147 -4079
rect -3141 -4083 -3137 -4079
rect -3124 -4083 -3120 -4079
rect -2547 -4048 -2543 -4044
rect -2530 -4048 -2526 -4044
rect -3106 -4153 -3102 -4149
rect -3089 -4153 -3085 -4149
rect -3113 -4527 -3109 -4523
rect -3057 -4514 -3053 -4510
rect -3040 -4514 -3036 -4510
rect -3113 -4544 -3109 -4540
rect -2996 -4526 -2992 -4522
rect -2979 -4526 -2975 -4522
rect -2969 -4526 -2965 -4522
rect -2952 -4526 -2948 -4522
rect -3113 -4578 -3109 -4574
rect -3113 -4595 -3109 -4591
rect -2934 -4596 -2930 -4592
rect -2917 -4596 -2913 -4592
rect -3165 -4706 -3161 -4702
rect -3148 -4706 -3144 -4702
rect -3138 -4706 -3134 -4702
rect -3121 -4706 -3117 -4702
rect -2848 -4730 -2844 -4726
rect -2831 -4730 -2827 -4726
rect -3103 -4776 -3099 -4772
rect -3086 -4776 -3082 -4772
rect -2799 -4778 -2795 -4774
rect -2782 -4778 -2778 -4774
<< polysilicon >>
rect 1785 412 1787 416
rect 1812 412 1814 416
rect 1785 367 1787 392
rect 1812 376 1814 392
rect 1804 338 1806 365
rect 1847 362 1849 365
rect 2143 342 2227 344
rect 1804 314 1806 318
rect 1847 295 1849 322
rect 2117 319 2120 321
rect 2130 319 2158 321
rect 2178 319 2183 321
rect 2225 317 2227 342
rect 2261 330 2263 336
rect 2225 304 2227 307
rect 2143 297 2227 299
rect 1804 283 1806 292
rect 2225 284 2227 297
rect 2261 292 2263 310
rect 1847 281 1849 284
rect 2261 275 2263 282
rect 2225 271 2227 274
rect 2117 268 2120 270
rect 2130 268 2158 270
rect 2178 268 2183 270
rect 2415 264 2417 274
rect 1804 260 1806 263
rect 2415 238 2417 244
rect 2415 236 2435 238
rect 2415 216 2417 225
rect 2415 191 2417 197
rect 2400 189 2417 191
rect 2400 172 2402 189
rect 2433 172 2435 236
rect 2464 220 2466 226
rect 2464 182 2466 200
rect 2464 165 2466 172
rect 2400 158 2402 162
rect 2433 158 2435 162
rect -3149 -2131 -3065 -2129
rect -3175 -2154 -3172 -2152
rect -3162 -2154 -3134 -2152
rect -3114 -2154 -3109 -2152
rect -3067 -2158 -3065 -2131
rect -3031 -2143 -3029 -2137
rect -3067 -2169 -3065 -2166
rect -3149 -2176 -3065 -2174
rect -3067 -2189 -3065 -2176
rect -3031 -2181 -3029 -2163
rect -2927 -2185 -2925 -2181
rect -2900 -2185 -2898 -2181
rect -3031 -2198 -3029 -2191
rect -3067 -2202 -3065 -2199
rect -3175 -2205 -3172 -2203
rect -3162 -2205 -3134 -2203
rect -3114 -2205 -3109 -2203
rect -2927 -2230 -2925 -2205
rect -2900 -2221 -2898 -2205
rect -2782 -2223 -2780 -2219
rect -2755 -2223 -2753 -2219
rect -2908 -2259 -2906 -2232
rect -2865 -2235 -2863 -2232
rect -2589 -2239 -2587 -2235
rect -2562 -2239 -2560 -2235
rect -2443 -2237 -2441 -2233
rect -2416 -2237 -2414 -2233
rect -2782 -2268 -2780 -2243
rect -2755 -2259 -2753 -2243
rect -2299 -2241 -2297 -2237
rect -2272 -2241 -2270 -2237
rect -2908 -2283 -2906 -2279
rect -2865 -2302 -2863 -2275
rect -2763 -2297 -2761 -2270
rect -2720 -2273 -2718 -2270
rect -2908 -2314 -2906 -2305
rect -2865 -2316 -2863 -2313
rect -2589 -2284 -2587 -2259
rect -2562 -2275 -2560 -2259
rect -2443 -2282 -2441 -2257
rect -2416 -2273 -2414 -2257
rect -2144 -2243 -2142 -2239
rect -2117 -2243 -2115 -2239
rect -2570 -2313 -2568 -2286
rect -2527 -2289 -2525 -2286
rect -2763 -2321 -2761 -2317
rect -2908 -2337 -2906 -2334
rect -2720 -2340 -2718 -2313
rect -2424 -2311 -2422 -2284
rect -2381 -2287 -2379 -2284
rect -2299 -2286 -2297 -2261
rect -2272 -2277 -2270 -2261
rect -2009 -2251 -2007 -2247
rect -1982 -2251 -1980 -2247
rect -2570 -2337 -2568 -2333
rect -3145 -2346 -3143 -2342
rect -3118 -2346 -3116 -2342
rect -2763 -2352 -2761 -2343
rect -3145 -2391 -3143 -2366
rect -3118 -2382 -3116 -2366
rect -2720 -2354 -2718 -2351
rect -2527 -2356 -2525 -2329
rect -2144 -2288 -2142 -2263
rect -2117 -2279 -2115 -2263
rect -2280 -2315 -2278 -2288
rect -2237 -2291 -2235 -2288
rect -2424 -2335 -2422 -2331
rect -2381 -2354 -2379 -2327
rect -2125 -2317 -2123 -2290
rect -2082 -2293 -2080 -2290
rect -2280 -2339 -2278 -2335
rect -2570 -2368 -2568 -2359
rect -2424 -2366 -2422 -2357
rect -2237 -2358 -2235 -2331
rect -2009 -2296 -2007 -2271
rect -1982 -2287 -1980 -2271
rect -1848 -2294 -1846 -2284
rect -1990 -2325 -1988 -2298
rect -1947 -2301 -1945 -2298
rect -2125 -2341 -2123 -2337
rect -2763 -2375 -2761 -2372
rect -2527 -2370 -2525 -2367
rect -2381 -2368 -2379 -2365
rect -2280 -2370 -2278 -2361
rect -2082 -2360 -2080 -2333
rect -1848 -2320 -1846 -2314
rect -1848 -2322 -1828 -2320
rect -1990 -2349 -1988 -2345
rect -2570 -2391 -2568 -2388
rect -2424 -2389 -2422 -2386
rect -2237 -2372 -2235 -2369
rect -2125 -2372 -2123 -2363
rect -1947 -2368 -1945 -2341
rect -1848 -2342 -1846 -2333
rect -1848 -2367 -1846 -2361
rect -2280 -2393 -2278 -2390
rect -2082 -2374 -2080 -2371
rect -1990 -2380 -1988 -2371
rect -1863 -2369 -1846 -2367
rect -3126 -2420 -3124 -2393
rect -3083 -2396 -3081 -2393
rect -2125 -2395 -2123 -2392
rect -1947 -2382 -1945 -2379
rect -1863 -2386 -1861 -2369
rect -1830 -2386 -1828 -2322
rect -1799 -2338 -1797 -2332
rect -1686 -2350 -1684 -2340
rect -1799 -2376 -1797 -2358
rect -1686 -2376 -1684 -2370
rect -1686 -2378 -1666 -2376
rect -1799 -2393 -1797 -2386
rect -1863 -2400 -1861 -2396
rect -1830 -2400 -1828 -2396
rect -1990 -2403 -1988 -2400
rect -1686 -2398 -1684 -2389
rect -1686 -2423 -1684 -2417
rect -1701 -2425 -1684 -2423
rect -3126 -2444 -3124 -2440
rect -3083 -2463 -3081 -2436
rect -1701 -2442 -1699 -2425
rect -1668 -2442 -1666 -2378
rect -1637 -2394 -1635 -2388
rect -1528 -2406 -1526 -2396
rect -1637 -2432 -1635 -2414
rect -1528 -2432 -1526 -2426
rect -1528 -2434 -1508 -2432
rect -1637 -2449 -1635 -2442
rect -1701 -2456 -1699 -2452
rect -1668 -2456 -1666 -2452
rect -1528 -2454 -1526 -2445
rect -3126 -2475 -3124 -2466
rect -3083 -2477 -3081 -2474
rect -1528 -2479 -1526 -2473
rect -1543 -2481 -1526 -2479
rect -3126 -2498 -3124 -2495
rect -1543 -2498 -1541 -2481
rect -1510 -2498 -1508 -2434
rect -1479 -2450 -1477 -2444
rect -1479 -2488 -1477 -2470
rect -1362 -2482 -1360 -2472
rect -1479 -2505 -1477 -2498
rect -1543 -2512 -1541 -2508
rect -1510 -2512 -1508 -2508
rect -1362 -2508 -1360 -2502
rect -1362 -2510 -1342 -2508
rect -1362 -2530 -1360 -2521
rect -1362 -2555 -1360 -2549
rect -1377 -2557 -1360 -2555
rect -1377 -2574 -1375 -2557
rect -1344 -2574 -1342 -2510
rect -1313 -2526 -1311 -2520
rect -1313 -2564 -1311 -2546
rect -1313 -2581 -1311 -2574
rect -1377 -2588 -1375 -2584
rect -1344 -2588 -1342 -2584
rect -3143 -2982 -3059 -2980
rect -3169 -3005 -3166 -3003
rect -3156 -3005 -3128 -3003
rect -3108 -3005 -3103 -3003
rect -3061 -3009 -3059 -2982
rect -3025 -2994 -3023 -2988
rect -2919 -3000 -2917 -2996
rect -2892 -3000 -2890 -2996
rect -2750 -2999 -2748 -2995
rect -2723 -2999 -2721 -2995
rect -2586 -2997 -2584 -2993
rect -2559 -2997 -2557 -2993
rect -3061 -3020 -3059 -3017
rect -3143 -3027 -3059 -3025
rect -3061 -3040 -3059 -3027
rect -3025 -3032 -3023 -3014
rect -2446 -2999 -2444 -2995
rect -2419 -2999 -2417 -2995
rect -3025 -3049 -3023 -3042
rect -2919 -3045 -2917 -3020
rect -2892 -3036 -2890 -3020
rect -2750 -3044 -2748 -3019
rect -2723 -3035 -2721 -3019
rect -2586 -3042 -2584 -3017
rect -2559 -3033 -2557 -3017
rect -2295 -3012 -2293 -3008
rect -2268 -3012 -2266 -3008
rect -2446 -3044 -2444 -3019
rect -2419 -3035 -2417 -3019
rect -3061 -3053 -3059 -3050
rect -3169 -3056 -3166 -3054
rect -3156 -3056 -3128 -3054
rect -3108 -3056 -3103 -3054
rect -2900 -3074 -2898 -3047
rect -2857 -3050 -2855 -3047
rect -2731 -3073 -2729 -3046
rect -2688 -3049 -2686 -3046
rect -2900 -3098 -2898 -3094
rect -2857 -3117 -2855 -3090
rect -2567 -3071 -2565 -3044
rect -2524 -3047 -2522 -3044
rect -2731 -3097 -2729 -3093
rect -2688 -3116 -2686 -3089
rect -2427 -3073 -2425 -3046
rect -2384 -3049 -2382 -3046
rect -2567 -3095 -2565 -3091
rect -2524 -3114 -2522 -3087
rect -2295 -3057 -2293 -3032
rect -2268 -3048 -2266 -3032
rect -1985 -3041 -1983 -3031
rect -2276 -3086 -2274 -3059
rect -2233 -3062 -2231 -3059
rect -2427 -3097 -2425 -3093
rect -2900 -3129 -2898 -3120
rect -2731 -3128 -2729 -3119
rect -2567 -3126 -2565 -3117
rect -2384 -3116 -2382 -3089
rect -1985 -3067 -1983 -3061
rect -1985 -3069 -1965 -3067
rect -1985 -3089 -1983 -3080
rect -2276 -3110 -2274 -3106
rect -2857 -3131 -2855 -3128
rect -2688 -3130 -2686 -3127
rect -2524 -3128 -2522 -3125
rect -2427 -3128 -2425 -3119
rect -2900 -3152 -2898 -3149
rect -2731 -3151 -2729 -3148
rect -2567 -3149 -2565 -3146
rect -2384 -3130 -2382 -3127
rect -2233 -3129 -2231 -3102
rect -1985 -3114 -1983 -3108
rect -2000 -3116 -1983 -3114
rect -2276 -3141 -2274 -3132
rect -2000 -3133 -1998 -3116
rect -1967 -3133 -1965 -3069
rect -1936 -3085 -1934 -3079
rect -1936 -3123 -1934 -3105
rect -2427 -3151 -2425 -3148
rect -2233 -3143 -2231 -3140
rect -1936 -3140 -1934 -3133
rect -2000 -3147 -1998 -3143
rect -1967 -3147 -1965 -3143
rect -2276 -3164 -2274 -3161
rect -2132 -3216 -2130 -3212
rect -2105 -3216 -2103 -3212
rect -3152 -3261 -3150 -3257
rect -3125 -3261 -3123 -3257
rect -2132 -3261 -2130 -3236
rect -2105 -3252 -2103 -3236
rect -1851 -3251 -1849 -3241
rect -3152 -3306 -3150 -3281
rect -3125 -3297 -3123 -3281
rect -2113 -3290 -2111 -3263
rect -2070 -3266 -2068 -3263
rect -3133 -3335 -3131 -3308
rect -3090 -3311 -3088 -3308
rect -1851 -3277 -1849 -3271
rect -1851 -3279 -1831 -3277
rect -1851 -3299 -1849 -3290
rect -2113 -3314 -2111 -3310
rect -2070 -3333 -2068 -3306
rect -1851 -3324 -1849 -3318
rect -1866 -3326 -1849 -3324
rect -2113 -3345 -2111 -3336
rect -1866 -3343 -1864 -3326
rect -1833 -3343 -1831 -3279
rect -1802 -3295 -1800 -3289
rect -1802 -3333 -1800 -3315
rect -3133 -3359 -3131 -3355
rect -3090 -3378 -3088 -3351
rect -2070 -3347 -2068 -3344
rect -1802 -3350 -1800 -3343
rect -1866 -3357 -1864 -3353
rect -1833 -3357 -1831 -3353
rect -2113 -3368 -2111 -3365
rect -3133 -3390 -3131 -3381
rect -3090 -3392 -3088 -3389
rect -3133 -3413 -3131 -3410
rect -1704 -3411 -1702 -3401
rect -1494 -3424 -1492 -3420
rect -1704 -3437 -1702 -3431
rect -1704 -3439 -1684 -3437
rect -1704 -3459 -1702 -3450
rect -1704 -3484 -1702 -3478
rect -1719 -3486 -1702 -3484
rect -1719 -3503 -1717 -3486
rect -1686 -3503 -1684 -3439
rect -1655 -3455 -1653 -3449
rect -1494 -3457 -1492 -3444
rect -1494 -3471 -1492 -3467
rect -1655 -3493 -1653 -3475
rect -1494 -3479 -1492 -3475
rect -1476 -3479 -1474 -3467
rect -1655 -3510 -1653 -3503
rect -1494 -3511 -1492 -3499
rect -1476 -3502 -1474 -3499
rect -1476 -3511 -1474 -3508
rect -1719 -3517 -1717 -3513
rect -1686 -3517 -1684 -3513
rect -1494 -3524 -1492 -3521
rect -1476 -3527 -1474 -3521
rect -3143 -3750 -3059 -3748
rect -3169 -3773 -3166 -3771
rect -3156 -3773 -3128 -3771
rect -3108 -3773 -3103 -3771
rect -3061 -3777 -3059 -3750
rect -3025 -3762 -3023 -3756
rect -2898 -3773 -2896 -3769
rect -2871 -3773 -2869 -3769
rect -3061 -3788 -3059 -3785
rect -3143 -3795 -3059 -3793
rect -3061 -3808 -3059 -3795
rect -3025 -3800 -3023 -3782
rect -3025 -3817 -3023 -3810
rect -2898 -3818 -2896 -3793
rect -2871 -3809 -2869 -3793
rect -3061 -3821 -3059 -3818
rect -3169 -3824 -3166 -3822
rect -3156 -3824 -3128 -3822
rect -3108 -3824 -3103 -3822
rect -2879 -3847 -2877 -3820
rect -2836 -3823 -2834 -3820
rect -2879 -3871 -2877 -3867
rect -2836 -3890 -2834 -3863
rect -2879 -3902 -2877 -3893
rect -2732 -3901 -2730 -3891
rect -2836 -3904 -2834 -3901
rect -2879 -3925 -2877 -3922
rect -2732 -3927 -2730 -3921
rect -2732 -3929 -2712 -3927
rect -2732 -3949 -2730 -3940
rect -2732 -3974 -2730 -3968
rect -2897 -3978 -2895 -3974
rect -2870 -3978 -2868 -3974
rect -2747 -3976 -2730 -3974
rect -2747 -3993 -2745 -3976
rect -2714 -3993 -2712 -3929
rect -2683 -3945 -2681 -3939
rect -2683 -3983 -2681 -3965
rect -2897 -4023 -2895 -3998
rect -2870 -4014 -2868 -3998
rect -2683 -4000 -2681 -3993
rect -2747 -4007 -2745 -4003
rect -2714 -4007 -2712 -4003
rect -2586 -4014 -2584 -4004
rect -2878 -4052 -2876 -4025
rect -2835 -4028 -2833 -4025
rect -2586 -4040 -2584 -4034
rect -2412 -4035 -2410 -4031
rect -2586 -4042 -2566 -4040
rect -2586 -4062 -2584 -4053
rect -2878 -4076 -2876 -4072
rect -2835 -4095 -2833 -4068
rect -2586 -4087 -2584 -4081
rect -2601 -4089 -2584 -4087
rect -3158 -4110 -3156 -4106
rect -3131 -4110 -3129 -4106
rect -2878 -4107 -2876 -4098
rect -2601 -4106 -2599 -4089
rect -2568 -4106 -2566 -4042
rect -2537 -4058 -2535 -4052
rect -2412 -4068 -2410 -4055
rect -2537 -4096 -2535 -4078
rect -2412 -4082 -2410 -4078
rect -2412 -4090 -2410 -4086
rect -2394 -4090 -2392 -4078
rect -2835 -4109 -2833 -4106
rect -2537 -4113 -2535 -4106
rect -2601 -4120 -2599 -4116
rect -2568 -4120 -2566 -4116
rect -2412 -4122 -2410 -4110
rect -2394 -4113 -2392 -4110
rect -2394 -4122 -2392 -4119
rect -2878 -4130 -2876 -4127
rect -3158 -4155 -3156 -4130
rect -3131 -4146 -3129 -4130
rect -2412 -4135 -2410 -4132
rect -2394 -4138 -2392 -4132
rect 713 -4135 715 -4131
rect -3139 -4184 -3137 -4157
rect -3096 -4160 -3094 -4157
rect 713 -4168 715 -4155
rect 713 -4182 715 -4178
rect 713 -4190 715 -4186
rect 731 -4190 733 -4178
rect -3139 -4208 -3137 -4204
rect -3096 -4227 -3094 -4200
rect 713 -4222 715 -4210
rect 731 -4213 733 -4210
rect 731 -4222 733 -4219
rect -3139 -4239 -3137 -4230
rect 713 -4235 715 -4232
rect 731 -4238 733 -4232
rect -3096 -4241 -3094 -4238
rect -3139 -4262 -3137 -4259
rect -3165 -4512 -3081 -4510
rect -3191 -4535 -3188 -4533
rect -3178 -4535 -3150 -4533
rect -3130 -4535 -3125 -4533
rect -3083 -4539 -3081 -4512
rect -3047 -4524 -3045 -4518
rect -3083 -4550 -3081 -4547
rect -3165 -4557 -3081 -4555
rect -3083 -4570 -3081 -4557
rect -3047 -4562 -3045 -4544
rect -2986 -4553 -2984 -4549
rect -2959 -4553 -2957 -4549
rect -3047 -4579 -3045 -4572
rect -3083 -4583 -3081 -4580
rect -3191 -4586 -3188 -4584
rect -3178 -4586 -3150 -4584
rect -3130 -4586 -3125 -4584
rect -2986 -4598 -2984 -4573
rect -2959 -4589 -2957 -4573
rect -2967 -4627 -2965 -4600
rect -2924 -4603 -2922 -4600
rect -2967 -4651 -2965 -4647
rect -2924 -4670 -2922 -4643
rect -2967 -4682 -2965 -4673
rect -2924 -4684 -2922 -4681
rect -2967 -4705 -2965 -4702
rect -3155 -4733 -3153 -4729
rect -3128 -4733 -3126 -4729
rect -2838 -4744 -2836 -4734
rect -3155 -4778 -3153 -4753
rect -3128 -4769 -3126 -4753
rect -2604 -4759 -2602 -4755
rect -2838 -4770 -2836 -4764
rect -2838 -4772 -2818 -4770
rect -3136 -4807 -3134 -4780
rect -3093 -4783 -3091 -4780
rect -2838 -4792 -2836 -4783
rect -2838 -4817 -2836 -4811
rect -2853 -4819 -2836 -4817
rect -3136 -4831 -3134 -4827
rect -3093 -4850 -3091 -4823
rect -2853 -4836 -2851 -4819
rect -2820 -4836 -2818 -4772
rect -2789 -4788 -2787 -4782
rect -2604 -4792 -2602 -4779
rect -2604 -4806 -2602 -4802
rect -2789 -4826 -2787 -4808
rect -2604 -4814 -2602 -4810
rect -2586 -4814 -2584 -4802
rect -2789 -4843 -2787 -4836
rect -2604 -4846 -2602 -4834
rect -2586 -4837 -2584 -4834
rect -2586 -4846 -2584 -4843
rect -2853 -4850 -2851 -4846
rect -2820 -4850 -2818 -4846
rect -3136 -4862 -3134 -4853
rect -2604 -4859 -2602 -4856
rect -3093 -4864 -3091 -4861
rect -2586 -4862 -2584 -4856
rect -2932 -4875 -2930 -4871
rect -3136 -4885 -3134 -4882
rect -2932 -4908 -2930 -4895
rect -2932 -4922 -2930 -4918
rect -2932 -4930 -2930 -4926
rect -2914 -4930 -2912 -4918
rect -2932 -4962 -2930 -4950
rect -2914 -4953 -2912 -4950
rect -2914 -4962 -2912 -4959
rect -2932 -4975 -2930 -4972
rect -2914 -4978 -2912 -4972
<< polycontact >>
rect 1780 370 1785 375
rect 1814 376 1819 380
rect 1798 360 1804 365
rect 2143 337 2148 342
rect 1842 307 1847 312
rect 2143 321 2148 326
rect 2143 299 2148 304
rect 1797 286 1804 291
rect 2256 295 2261 300
rect 2143 270 2148 275
rect 2410 236 2415 241
rect 2395 186 2400 191
rect 2459 185 2464 190
rect -3149 -2136 -3144 -2131
rect -3149 -2152 -3144 -2147
rect -3149 -2174 -3144 -2169
rect -3036 -2178 -3031 -2173
rect -3149 -2203 -3144 -2198
rect -2932 -2227 -2927 -2222
rect -2898 -2221 -2893 -2217
rect -2914 -2237 -2908 -2232
rect -2787 -2265 -2782 -2260
rect -2753 -2259 -2748 -2255
rect -2769 -2275 -2763 -2270
rect -2870 -2290 -2865 -2285
rect -2915 -2311 -2908 -2306
rect -2594 -2281 -2589 -2276
rect -2560 -2275 -2555 -2271
rect -2448 -2279 -2443 -2274
rect -2414 -2273 -2409 -2269
rect -2304 -2283 -2299 -2278
rect -2576 -2291 -2570 -2286
rect -2430 -2289 -2424 -2284
rect -2725 -2328 -2720 -2323
rect -2270 -2277 -2265 -2273
rect -2149 -2285 -2144 -2280
rect -2770 -2349 -2763 -2344
rect -2532 -2344 -2527 -2339
rect -3150 -2388 -3145 -2383
rect -2115 -2279 -2110 -2275
rect -2286 -2293 -2280 -2288
rect -2386 -2342 -2381 -2337
rect -2131 -2295 -2125 -2290
rect -2014 -2293 -2009 -2288
rect -2242 -2346 -2237 -2341
rect -2577 -2365 -2570 -2360
rect -2431 -2363 -2424 -2358
rect -1980 -2287 -1975 -2283
rect -1996 -2303 -1990 -2298
rect -2087 -2348 -2082 -2343
rect -3116 -2382 -3111 -2378
rect -2287 -2367 -2280 -2362
rect -1853 -2322 -1848 -2317
rect -1952 -2356 -1947 -2351
rect -2132 -2369 -2125 -2364
rect -1997 -2377 -1990 -2372
rect -1868 -2372 -1863 -2367
rect -3132 -2398 -3126 -2393
rect -1804 -2373 -1799 -2368
rect -1691 -2378 -1686 -2373
rect -1706 -2428 -1701 -2423
rect -3088 -2451 -3083 -2446
rect -1642 -2429 -1637 -2424
rect -1533 -2434 -1528 -2429
rect -3133 -2472 -3126 -2467
rect -1548 -2484 -1543 -2479
rect -1484 -2485 -1479 -2480
rect -1367 -2510 -1362 -2505
rect -1382 -2560 -1377 -2555
rect -1318 -2561 -1313 -2556
rect -3143 -2987 -3138 -2982
rect -3143 -3003 -3138 -2998
rect -3143 -3025 -3138 -3020
rect -3030 -3029 -3025 -3024
rect -3143 -3054 -3138 -3049
rect -2924 -3042 -2919 -3037
rect -2890 -3036 -2885 -3032
rect -2755 -3041 -2750 -3036
rect -2721 -3035 -2716 -3031
rect -2591 -3039 -2586 -3034
rect -2557 -3033 -2552 -3029
rect -2451 -3041 -2446 -3036
rect -2417 -3035 -2412 -3031
rect -2906 -3052 -2900 -3047
rect -2737 -3051 -2731 -3046
rect -2573 -3049 -2567 -3044
rect -2862 -3105 -2857 -3100
rect -2693 -3104 -2688 -3099
rect -2433 -3051 -2427 -3046
rect -2529 -3102 -2524 -3097
rect -2300 -3054 -2295 -3049
rect -2266 -3048 -2261 -3044
rect -2282 -3064 -2276 -3059
rect -2389 -3104 -2384 -3099
rect -2907 -3126 -2900 -3121
rect -2738 -3125 -2731 -3120
rect -2574 -3123 -2567 -3118
rect -1990 -3069 -1985 -3064
rect -2434 -3125 -2427 -3120
rect -2238 -3117 -2233 -3112
rect -2005 -3119 -2000 -3114
rect -2283 -3138 -2276 -3133
rect -1941 -3120 -1936 -3115
rect -2137 -3258 -2132 -3253
rect -2103 -3252 -2098 -3248
rect -2119 -3268 -2113 -3263
rect -3157 -3303 -3152 -3298
rect -3123 -3297 -3118 -3293
rect -3139 -3313 -3133 -3308
rect -1856 -3279 -1851 -3274
rect -2075 -3321 -2070 -3316
rect -1871 -3329 -1866 -3324
rect -2120 -3342 -2113 -3337
rect -1807 -3330 -1802 -3325
rect -3095 -3366 -3090 -3361
rect -3140 -3387 -3133 -3382
rect -1709 -3439 -1704 -3434
rect -1724 -3489 -1719 -3484
rect -1498 -3456 -1494 -3452
rect -1480 -3472 -1476 -3468
rect -1660 -3490 -1655 -3485
rect -1498 -3510 -1494 -3506
rect -1474 -3526 -1470 -3522
rect -3143 -3755 -3138 -3750
rect -3143 -3771 -3138 -3766
rect -3143 -3793 -3138 -3788
rect -3030 -3797 -3025 -3792
rect -3143 -3822 -3138 -3817
rect -2903 -3815 -2898 -3810
rect -2869 -3809 -2864 -3805
rect -2885 -3825 -2879 -3820
rect -2841 -3878 -2836 -3873
rect -2886 -3899 -2879 -3894
rect -2737 -3929 -2732 -3924
rect -2752 -3979 -2747 -3974
rect -2688 -3980 -2683 -3975
rect -2902 -4020 -2897 -4015
rect -2868 -4014 -2863 -4010
rect -2884 -4030 -2878 -4025
rect -2591 -4042 -2586 -4037
rect -2840 -4083 -2835 -4078
rect -2606 -4092 -2601 -4087
rect -2885 -4104 -2878 -4099
rect -2416 -4067 -2412 -4063
rect -2542 -4093 -2537 -4088
rect -2398 -4083 -2394 -4079
rect -2416 -4121 -2412 -4117
rect -3163 -4152 -3158 -4147
rect -2392 -4137 -2388 -4133
rect -3129 -4146 -3124 -4142
rect -3145 -4162 -3139 -4157
rect 709 -4167 713 -4163
rect 727 -4183 731 -4179
rect -3101 -4215 -3096 -4210
rect 709 -4221 713 -4217
rect -3146 -4236 -3139 -4231
rect 733 -4237 737 -4233
rect -3165 -4517 -3160 -4512
rect -3165 -4533 -3160 -4528
rect -3165 -4555 -3160 -4550
rect -3052 -4559 -3047 -4554
rect -3165 -4584 -3160 -4579
rect -2991 -4595 -2986 -4590
rect -2957 -4589 -2952 -4585
rect -2973 -4605 -2967 -4600
rect -2929 -4658 -2924 -4653
rect -2974 -4679 -2967 -4674
rect -3160 -4775 -3155 -4770
rect -3126 -4769 -3121 -4765
rect -2843 -4772 -2838 -4767
rect -3142 -4785 -3136 -4780
rect -2858 -4822 -2853 -4817
rect -3098 -4838 -3093 -4833
rect -2608 -4791 -2604 -4787
rect -2590 -4807 -2586 -4803
rect -2794 -4823 -2789 -4818
rect -2608 -4845 -2604 -4841
rect -3143 -4859 -3136 -4854
rect -2584 -4861 -2580 -4857
rect -2936 -4907 -2932 -4903
rect -2918 -4923 -2914 -4919
rect -2936 -4961 -2932 -4957
rect -2912 -4977 -2908 -4973
<< metal1 >>
rect 1772 443 1826 446
rect 1772 439 1775 443
rect 1779 439 1792 443
rect 1796 439 1802 443
rect 1806 439 1819 443
rect 1823 439 1826 443
rect 1772 437 1826 439
rect 1780 412 1784 437
rect 1815 412 1819 437
rect 1767 370 1780 375
rect 1788 372 1792 392
rect 1807 372 1811 392
rect 1819 376 1826 380
rect 1767 365 1772 370
rect 1788 368 1811 372
rect 1821 368 1826 376
rect 1834 373 1861 376
rect 1834 369 1837 373
rect 1841 369 1854 373
rect 1858 369 1861 373
rect 1767 360 1798 365
rect 1767 347 1772 360
rect 1759 344 1772 347
rect 1807 348 1811 368
rect 1834 367 1861 369
rect 1842 362 1846 367
rect 1807 342 1830 348
rect 1807 338 1811 342
rect 1799 312 1803 318
rect 1824 312 1830 342
rect 2248 344 2275 347
rect 2117 337 2143 342
rect 2248 340 2251 344
rect 2255 340 2268 344
rect 2272 340 2275 344
rect 2248 338 2275 340
rect 1850 312 1854 322
rect 2108 333 2114 334
rect 2108 329 2109 333
rect 2113 329 2114 333
rect 2108 326 2114 329
rect 2143 326 2148 337
rect 2193 331 2202 334
rect 2193 327 2195 331
rect 2199 327 2202 331
rect 2193 326 2202 327
rect 2108 322 2120 326
rect 2108 312 2114 322
rect 2178 322 2202 326
rect 2256 330 2260 338
rect 2143 314 2158 318
rect 2193 314 2202 322
rect 2228 318 2241 322
rect 2228 317 2232 318
rect 1799 308 1811 312
rect 1772 291 1778 292
rect 1772 286 1785 291
rect 1791 286 1797 291
rect 1807 283 1811 308
rect 1824 307 1842 312
rect 1850 307 1863 312
rect 2108 308 2109 312
rect 2113 308 2114 312
rect 2108 307 2114 308
rect 1850 295 1854 307
rect 2143 304 2148 314
rect 2193 310 2195 314
rect 2199 310 2202 314
rect 2193 307 2202 310
rect 2220 304 2224 307
rect 2172 300 2224 304
rect 2172 295 2176 300
rect 2113 290 2176 295
rect 1842 278 1846 284
rect 2108 282 2114 283
rect 2108 278 2109 282
rect 2113 278 2114 282
rect 1834 277 1861 278
rect 1834 273 1835 277
rect 1839 273 1856 277
rect 1860 273 1861 277
rect 1834 272 1861 273
rect 2108 275 2114 278
rect 2143 275 2148 290
rect 2228 284 2232 307
rect 2235 300 2241 318
rect 2264 300 2268 310
rect 2235 295 2256 300
rect 2264 295 2274 300
rect 2264 292 2268 295
rect 2193 280 2202 283
rect 2193 276 2195 280
rect 2199 276 2202 280
rect 2193 275 2202 276
rect 2108 271 2120 275
rect 1799 257 1803 263
rect 2108 261 2114 271
rect 2178 271 2202 275
rect 2143 263 2158 267
rect 2193 263 2202 271
rect 2108 257 2109 261
rect 2113 257 2114 261
rect 1791 256 1818 257
rect 2108 256 2114 257
rect 1791 252 1792 256
rect 1796 252 1813 256
rect 1817 252 1818 256
rect 1791 251 1818 252
rect 2143 252 2148 263
rect 2193 259 2195 263
rect 2199 259 2202 263
rect 2193 256 2202 259
rect 2402 282 2429 285
rect 2220 252 2224 274
rect 2256 272 2260 282
rect 2402 278 2405 282
rect 2409 278 2422 282
rect 2426 278 2429 282
rect 2402 276 2429 278
rect 2248 271 2275 272
rect 2248 267 2249 271
rect 2253 267 2270 271
rect 2274 267 2275 271
rect 2248 266 2275 267
rect 2143 249 2224 252
rect 2410 264 2414 276
rect 2393 236 2410 241
rect 2418 232 2422 244
rect 2410 228 2422 232
rect 2451 234 2478 237
rect 2451 230 2454 234
rect 2458 230 2471 234
rect 2475 230 2478 234
rect 2451 228 2478 230
rect 2410 216 2414 228
rect 2459 220 2463 228
rect 2386 186 2395 191
rect 2418 190 2422 197
rect 2467 190 2471 200
rect 2418 185 2459 190
rect 2467 185 2480 190
rect 2418 182 2422 185
rect 2467 182 2471 185
rect 2403 178 2440 182
rect 2403 172 2407 178
rect 2436 172 2440 178
rect 2459 162 2463 172
rect 2395 155 2399 162
rect 2428 155 2432 162
rect 2451 161 2478 162
rect 2451 157 2452 161
rect 2456 157 2473 161
rect 2477 157 2478 161
rect 2451 156 2478 157
rect 2387 154 2414 155
rect 2387 150 2388 154
rect 2392 150 2409 154
rect 2413 150 2414 154
rect 2387 149 2414 150
rect 2420 154 2447 155
rect 2420 150 2421 154
rect 2425 150 2442 154
rect 2446 150 2447 154
rect 2420 149 2447 150
rect -2987 -2108 -2970 -2103
rect -2961 -2108 -2040 -2103
rect -3044 -2129 -3017 -2126
rect -3262 -2136 -3149 -2131
rect -3044 -2133 -3041 -2129
rect -3037 -2133 -3024 -2129
rect -3020 -2133 -3017 -2129
rect -3044 -2135 -3017 -2133
rect -3262 -2409 -3257 -2136
rect -3184 -2140 -3178 -2139
rect -3184 -2144 -3183 -2140
rect -3179 -2144 -3178 -2140
rect -3184 -2147 -3178 -2144
rect -3149 -2147 -3144 -2136
rect -3099 -2142 -3090 -2139
rect -3099 -2146 -3097 -2142
rect -3093 -2146 -3090 -2142
rect -3099 -2147 -3090 -2146
rect -3184 -2151 -3172 -2147
rect -3184 -2161 -3178 -2151
rect -3114 -2151 -3090 -2147
rect -3036 -2143 -3032 -2135
rect -3149 -2159 -3134 -2155
rect -3099 -2159 -3090 -2151
rect -3064 -2155 -3051 -2151
rect -3064 -2158 -3060 -2155
rect -3184 -2165 -3183 -2161
rect -3179 -2165 -3178 -2161
rect -3184 -2166 -3178 -2165
rect -3149 -2169 -3144 -2159
rect -3099 -2163 -3097 -2159
rect -3093 -2163 -3090 -2159
rect -3099 -2166 -3090 -2163
rect -3072 -2169 -3068 -2166
rect -3120 -2173 -3068 -2169
rect -3120 -2178 -3116 -2173
rect -3175 -2183 -3116 -2178
rect -3184 -2191 -3178 -2190
rect -3184 -2195 -3183 -2191
rect -3179 -2195 -3178 -2191
rect -3184 -2198 -3178 -2195
rect -3149 -2198 -3144 -2183
rect -3064 -2189 -3060 -2166
rect -3057 -2173 -3051 -2155
rect -3028 -2173 -3024 -2163
rect -2987 -2173 -2982 -2108
rect -2940 -2154 -2886 -2151
rect -2940 -2158 -2937 -2154
rect -2933 -2158 -2920 -2154
rect -2916 -2158 -2910 -2154
rect -2906 -2158 -2893 -2154
rect -2889 -2158 -2886 -2154
rect -2940 -2160 -2886 -2158
rect -3057 -2178 -3036 -2173
rect -3028 -2178 -2982 -2173
rect -3028 -2181 -3024 -2178
rect -3099 -2193 -3090 -2190
rect -3099 -2197 -3097 -2193
rect -3093 -2197 -3090 -2193
rect -3099 -2198 -3090 -2197
rect -3184 -2202 -3172 -2198
rect -3184 -2212 -3178 -2202
rect -3114 -2202 -3090 -2198
rect -3149 -2210 -3134 -2206
rect -3099 -2210 -3090 -2202
rect -3184 -2216 -3183 -2212
rect -3179 -2216 -3178 -2212
rect -3184 -2217 -3178 -2216
rect -3149 -2221 -3144 -2210
rect -3099 -2214 -3097 -2210
rect -3093 -2214 -3090 -2210
rect -3099 -2217 -3090 -2214
rect -2932 -2185 -2928 -2160
rect -2897 -2185 -2893 -2160
rect -3072 -2221 -3068 -2199
rect -3036 -2201 -3032 -2191
rect -3044 -2202 -3017 -2201
rect -3044 -2206 -3043 -2202
rect -3039 -2206 -3022 -2202
rect -3018 -2206 -3017 -2202
rect -3044 -2207 -3017 -2206
rect -3149 -2224 -3068 -2221
rect -2945 -2227 -2932 -2222
rect -2924 -2225 -2920 -2205
rect -2905 -2225 -2901 -2205
rect -2893 -2221 -2886 -2217
rect -2945 -2232 -2940 -2227
rect -2924 -2229 -2901 -2225
rect -2891 -2229 -2886 -2221
rect -2878 -2224 -2851 -2221
rect -2878 -2228 -2875 -2224
rect -2871 -2228 -2858 -2224
rect -2854 -2228 -2851 -2224
rect -2945 -2237 -2914 -2232
rect -2945 -2248 -2940 -2237
rect -3006 -2253 -2940 -2248
rect -2905 -2249 -2901 -2229
rect -2878 -2230 -2851 -2228
rect -2870 -2235 -2866 -2230
rect -3158 -2315 -3104 -2312
rect -3158 -2319 -3155 -2315
rect -3151 -2319 -3138 -2315
rect -3134 -2319 -3128 -2315
rect -3124 -2319 -3111 -2315
rect -3107 -2319 -3104 -2315
rect -3158 -2321 -3104 -2319
rect -3150 -2346 -3146 -2321
rect -3115 -2346 -3111 -2321
rect -3163 -2388 -3150 -2383
rect -3142 -2386 -3138 -2366
rect -3123 -2386 -3119 -2366
rect -3111 -2382 -3104 -2378
rect -3163 -2393 -3158 -2388
rect -3142 -2390 -3119 -2386
rect -3109 -2390 -3104 -2382
rect -3096 -2385 -3069 -2382
rect -3096 -2389 -3093 -2385
rect -3089 -2389 -3076 -2385
rect -3072 -2389 -3069 -2385
rect -3163 -2398 -3132 -2393
rect -3163 -2409 -3158 -2398
rect -3262 -2414 -3158 -2409
rect -3123 -2410 -3119 -2390
rect -3096 -2391 -3069 -2389
rect -3088 -2396 -3084 -2391
rect -3123 -2416 -3100 -2410
rect -3123 -2420 -3119 -2416
rect -3131 -2446 -3127 -2440
rect -3106 -2446 -3100 -2416
rect -3080 -2446 -3076 -2436
rect -3131 -2450 -3119 -2446
rect -3158 -2451 -3152 -2450
rect -3158 -2467 -3152 -2456
rect -3158 -2472 -3145 -2467
rect -3139 -2472 -3133 -2467
rect -3123 -2475 -3119 -2450
rect -3106 -2451 -3088 -2446
rect -3080 -2451 -3073 -2446
rect -3080 -2463 -3076 -2451
rect -3088 -2480 -3084 -2474
rect -3096 -2481 -3069 -2480
rect -3096 -2485 -3095 -2481
rect -3091 -2485 -3074 -2481
rect -3070 -2485 -3069 -2481
rect -3096 -2486 -3069 -2485
rect -3131 -2501 -3127 -2495
rect -3139 -2502 -3112 -2501
rect -3139 -2506 -3138 -2502
rect -3134 -2506 -3117 -2502
rect -3113 -2506 -3112 -2502
rect -3139 -2507 -3112 -2506
rect -3006 -2917 -3001 -2253
rect -2905 -2255 -2882 -2249
rect -2905 -2259 -2901 -2255
rect -2913 -2285 -2909 -2279
rect -2888 -2285 -2882 -2255
rect -2862 -2285 -2858 -2275
rect -2913 -2289 -2901 -2285
rect -2974 -2306 -2934 -2305
rect -2974 -2309 -2927 -2306
rect -2974 -2867 -2970 -2309
rect -2940 -2311 -2927 -2309
rect -2921 -2311 -2915 -2306
rect -2905 -2314 -2901 -2289
rect -2888 -2290 -2870 -2285
rect -2862 -2290 -2832 -2285
rect -2862 -2302 -2858 -2290
rect -2870 -2319 -2866 -2313
rect -2878 -2320 -2851 -2319
rect -2878 -2324 -2877 -2320
rect -2873 -2324 -2856 -2320
rect -2852 -2324 -2851 -2320
rect -2878 -2325 -2851 -2324
rect -2913 -2340 -2909 -2334
rect -2921 -2341 -2894 -2340
rect -2921 -2345 -2920 -2341
rect -2916 -2345 -2899 -2341
rect -2895 -2345 -2894 -2341
rect -2921 -2346 -2894 -2345
rect -2837 -2343 -2832 -2290
rect -2819 -2287 -2814 -2108
rect -2795 -2192 -2741 -2189
rect -2795 -2196 -2792 -2192
rect -2788 -2196 -2775 -2192
rect -2771 -2196 -2765 -2192
rect -2761 -2196 -2748 -2192
rect -2744 -2196 -2741 -2192
rect -2795 -2198 -2741 -2196
rect -2787 -2223 -2783 -2198
rect -2752 -2223 -2748 -2198
rect -2602 -2208 -2548 -2205
rect -2602 -2212 -2599 -2208
rect -2595 -2212 -2582 -2208
rect -2578 -2212 -2572 -2208
rect -2568 -2212 -2555 -2208
rect -2551 -2212 -2548 -2208
rect -2602 -2214 -2548 -2212
rect -2800 -2265 -2787 -2260
rect -2779 -2263 -2775 -2243
rect -2594 -2239 -2590 -2214
rect -2559 -2239 -2555 -2214
rect -2760 -2263 -2756 -2243
rect -2748 -2259 -2741 -2255
rect -2800 -2270 -2795 -2265
rect -2779 -2267 -2756 -2263
rect -2746 -2267 -2741 -2259
rect -2733 -2262 -2706 -2259
rect -2733 -2266 -2730 -2262
rect -2726 -2266 -2713 -2262
rect -2709 -2266 -2706 -2262
rect -2800 -2275 -2769 -2270
rect -2800 -2287 -2795 -2275
rect -2819 -2292 -2795 -2287
rect -2760 -2287 -2756 -2267
rect -2733 -2268 -2706 -2266
rect -2725 -2273 -2721 -2268
rect -2760 -2293 -2737 -2287
rect -2760 -2297 -2756 -2293
rect -2768 -2323 -2764 -2317
rect -2743 -2323 -2737 -2293
rect -2607 -2281 -2594 -2276
rect -2586 -2279 -2582 -2259
rect -2567 -2279 -2563 -2259
rect -2555 -2275 -2548 -2271
rect -2607 -2286 -2602 -2281
rect -2586 -2283 -2563 -2279
rect -2553 -2283 -2548 -2275
rect -2540 -2278 -2513 -2275
rect -2540 -2282 -2537 -2278
rect -2533 -2282 -2520 -2278
rect -2516 -2282 -2513 -2278
rect -2607 -2291 -2576 -2286
rect -2607 -2303 -2602 -2291
rect -2717 -2323 -2713 -2313
rect -2682 -2308 -2602 -2303
rect -2567 -2303 -2563 -2283
rect -2540 -2284 -2513 -2282
rect -2532 -2289 -2528 -2284
rect -2768 -2327 -2756 -2323
rect -2837 -2344 -2787 -2343
rect -2837 -2349 -2782 -2344
rect -2776 -2349 -2770 -2344
rect -2837 -2351 -2787 -2349
rect -2760 -2352 -2756 -2327
rect -2743 -2328 -2725 -2323
rect -2717 -2328 -2710 -2323
rect -2717 -2340 -2713 -2328
rect -2725 -2357 -2721 -2351
rect -2733 -2358 -2706 -2357
rect -2733 -2362 -2732 -2358
rect -2728 -2362 -2711 -2358
rect -2707 -2362 -2706 -2358
rect -2733 -2363 -2706 -2362
rect -2768 -2378 -2764 -2372
rect -2776 -2379 -2749 -2378
rect -2776 -2383 -2775 -2379
rect -2771 -2383 -2754 -2379
rect -2750 -2383 -2749 -2379
rect -2776 -2384 -2749 -2383
rect -2682 -2727 -2677 -2308
rect -2634 -2410 -2629 -2308
rect -2567 -2309 -2544 -2303
rect -2567 -2313 -2563 -2309
rect -2575 -2339 -2571 -2333
rect -2550 -2339 -2544 -2309
rect -2486 -2300 -2481 -2108
rect -2456 -2206 -2402 -2203
rect -2456 -2210 -2453 -2206
rect -2449 -2210 -2436 -2206
rect -2432 -2210 -2426 -2206
rect -2422 -2210 -2409 -2206
rect -2405 -2210 -2402 -2206
rect -2456 -2212 -2402 -2210
rect -2312 -2210 -2258 -2207
rect -2448 -2237 -2444 -2212
rect -2413 -2237 -2409 -2212
rect -2312 -2214 -2309 -2210
rect -2305 -2214 -2292 -2210
rect -2288 -2214 -2282 -2210
rect -2278 -2214 -2265 -2210
rect -2261 -2214 -2258 -2210
rect -2312 -2216 -2258 -2214
rect -2461 -2279 -2448 -2274
rect -2440 -2277 -2436 -2257
rect -2304 -2241 -2300 -2216
rect -2269 -2241 -2265 -2216
rect -2421 -2277 -2417 -2257
rect -2409 -2273 -2402 -2269
rect -2461 -2284 -2456 -2279
rect -2440 -2281 -2417 -2277
rect -2407 -2281 -2402 -2273
rect -2394 -2276 -2367 -2273
rect -2394 -2280 -2391 -2276
rect -2387 -2280 -2374 -2276
rect -2370 -2280 -2367 -2276
rect -2461 -2289 -2430 -2284
rect -2461 -2300 -2456 -2289
rect -2486 -2305 -2456 -2300
rect -2421 -2301 -2417 -2281
rect -2394 -2282 -2367 -2280
rect -2386 -2287 -2382 -2282
rect -2317 -2283 -2304 -2278
rect -2296 -2281 -2292 -2261
rect -2277 -2281 -2273 -2261
rect -2265 -2277 -2258 -2273
rect -2421 -2307 -2398 -2301
rect -2421 -2311 -2417 -2307
rect -2524 -2339 -2520 -2329
rect -2429 -2337 -2425 -2331
rect -2404 -2337 -2398 -2307
rect -2317 -2288 -2312 -2283
rect -2296 -2285 -2273 -2281
rect -2263 -2285 -2258 -2277
rect -2250 -2280 -2223 -2277
rect -2250 -2284 -2247 -2280
rect -2243 -2284 -2230 -2280
rect -2226 -2284 -2223 -2280
rect -2317 -2293 -2286 -2288
rect -2317 -2311 -2312 -2293
rect -2277 -2305 -2273 -2285
rect -2250 -2286 -2223 -2284
rect -2242 -2291 -2238 -2286
rect -2277 -2311 -2254 -2305
rect -2277 -2315 -2273 -2311
rect -2378 -2337 -2374 -2327
rect -2575 -2343 -2563 -2339
rect -2594 -2365 -2589 -2360
rect -2583 -2365 -2577 -2360
rect -2567 -2368 -2563 -2343
rect -2550 -2344 -2532 -2339
rect -2524 -2344 -2450 -2339
rect -2429 -2341 -2417 -2337
rect -2524 -2356 -2520 -2344
rect -2455 -2358 -2450 -2344
rect -2455 -2363 -2443 -2358
rect -2437 -2363 -2431 -2358
rect -2421 -2366 -2417 -2341
rect -2404 -2342 -2386 -2337
rect -2378 -2342 -2326 -2337
rect -2378 -2354 -2374 -2342
rect -2532 -2373 -2528 -2367
rect -2540 -2374 -2513 -2373
rect -2540 -2378 -2539 -2374
rect -2535 -2378 -2518 -2374
rect -2514 -2378 -2513 -2374
rect -2540 -2379 -2513 -2378
rect -2386 -2371 -2382 -2365
rect -2394 -2372 -2367 -2371
rect -2394 -2376 -2393 -2372
rect -2389 -2376 -2372 -2372
rect -2368 -2376 -2367 -2372
rect -2394 -2377 -2367 -2376
rect -2575 -2394 -2571 -2388
rect -2429 -2392 -2425 -2386
rect -2437 -2393 -2410 -2392
rect -2583 -2395 -2556 -2394
rect -2583 -2399 -2582 -2395
rect -2578 -2399 -2561 -2395
rect -2557 -2399 -2556 -2395
rect -2437 -2397 -2436 -2393
rect -2432 -2397 -2415 -2393
rect -2411 -2397 -2410 -2393
rect -2437 -2398 -2410 -2397
rect -2331 -2393 -2326 -2342
rect -2285 -2341 -2281 -2335
rect -2260 -2341 -2254 -2311
rect -2200 -2307 -2195 -2108
rect -2157 -2212 -2103 -2209
rect -2157 -2216 -2154 -2212
rect -2150 -2216 -2137 -2212
rect -2133 -2216 -2127 -2212
rect -2123 -2216 -2110 -2212
rect -2106 -2216 -2103 -2212
rect -2157 -2218 -2103 -2216
rect -2149 -2243 -2145 -2218
rect -2114 -2243 -2110 -2218
rect -2162 -2285 -2149 -2280
rect -2141 -2283 -2137 -2263
rect -2122 -2283 -2118 -2263
rect -2110 -2279 -2103 -2275
rect -2162 -2290 -2157 -2285
rect -2141 -2287 -2118 -2283
rect -2108 -2287 -2103 -2279
rect -2095 -2282 -2068 -2279
rect -2095 -2286 -2092 -2282
rect -2088 -2286 -2075 -2282
rect -2071 -2286 -2068 -2282
rect -2162 -2295 -2131 -2290
rect -2162 -2307 -2157 -2295
rect -2200 -2312 -2157 -2307
rect -2122 -2307 -2118 -2287
rect -2095 -2288 -2068 -2286
rect -2087 -2293 -2083 -2288
rect -2122 -2313 -2099 -2307
rect -2122 -2317 -2118 -2313
rect -2234 -2341 -2230 -2331
rect -2285 -2345 -2273 -2341
rect -2313 -2362 -2306 -2361
rect -2313 -2367 -2299 -2362
rect -2293 -2367 -2287 -2362
rect -2583 -2400 -2556 -2399
rect -2313 -2410 -2308 -2367
rect -2277 -2370 -2273 -2345
rect -2260 -2346 -2242 -2341
rect -2234 -2346 -2188 -2341
rect -2234 -2358 -2230 -2346
rect -2193 -2363 -2188 -2346
rect -2130 -2343 -2126 -2337
rect -2105 -2343 -2099 -2313
rect -2045 -2314 -2040 -2108
rect -2022 -2220 -1968 -2217
rect -2022 -2224 -2019 -2220
rect -2015 -2224 -2002 -2220
rect -1998 -2224 -1992 -2220
rect -1988 -2224 -1975 -2220
rect -1971 -2224 -1968 -2220
rect -2022 -2226 -1968 -2224
rect -2014 -2251 -2010 -2226
rect -1979 -2251 -1975 -2226
rect -2027 -2293 -2014 -2288
rect -2006 -2291 -2002 -2271
rect -1889 -2249 -1569 -2244
rect -1987 -2291 -1983 -2271
rect -1975 -2287 -1968 -2283
rect -2027 -2298 -2022 -2293
rect -2006 -2295 -1983 -2291
rect -1973 -2295 -1968 -2287
rect -1960 -2290 -1933 -2287
rect -1960 -2294 -1957 -2290
rect -1953 -2294 -1940 -2290
rect -1936 -2294 -1933 -2290
rect -2027 -2303 -1996 -2298
rect -2027 -2314 -2022 -2303
rect -2045 -2319 -2021 -2314
rect -1987 -2315 -1983 -2295
rect -1960 -2296 -1933 -2294
rect -1952 -2301 -1948 -2296
rect -1987 -2321 -1964 -2315
rect -1987 -2325 -1983 -2321
rect -2079 -2343 -2075 -2333
rect -2130 -2347 -2118 -2343
rect -2193 -2364 -2145 -2363
rect -2193 -2368 -2144 -2364
rect -2157 -2369 -2144 -2368
rect -2138 -2369 -2132 -2364
rect -2242 -2375 -2238 -2369
rect -2122 -2372 -2118 -2347
rect -2105 -2348 -2087 -2343
rect -2079 -2348 -2041 -2343
rect -2079 -2360 -2075 -2348
rect -2250 -2376 -2223 -2375
rect -2250 -2380 -2249 -2376
rect -2245 -2380 -2228 -2376
rect -2224 -2380 -2223 -2376
rect -2250 -2381 -2223 -2380
rect -2285 -2396 -2281 -2390
rect -2087 -2377 -2083 -2371
rect -2095 -2378 -2068 -2377
rect -2095 -2382 -2094 -2378
rect -2090 -2382 -2073 -2378
rect -2069 -2382 -2068 -2378
rect -2095 -2383 -2068 -2382
rect -2293 -2397 -2266 -2396
rect -2293 -2401 -2292 -2397
rect -2288 -2401 -2271 -2397
rect -2267 -2401 -2266 -2397
rect -2130 -2398 -2126 -2392
rect -2293 -2402 -2266 -2401
rect -2138 -2399 -2111 -2398
rect -2138 -2403 -2137 -2399
rect -2133 -2403 -2116 -2399
rect -2112 -2403 -2111 -2399
rect -2138 -2404 -2111 -2403
rect -2634 -2415 -2308 -2410
rect -2046 -2447 -2041 -2348
rect -1995 -2351 -1991 -2345
rect -1970 -2351 -1964 -2321
rect -1944 -2351 -1940 -2341
rect -1889 -2351 -1884 -2249
rect -1861 -2276 -1834 -2273
rect -1861 -2280 -1858 -2276
rect -1854 -2280 -1841 -2276
rect -1837 -2280 -1834 -2276
rect -1861 -2282 -1834 -2280
rect -1853 -2294 -1849 -2282
rect -1864 -2322 -1853 -2317
rect -1845 -2326 -1841 -2314
rect -1995 -2355 -1983 -2351
rect -2022 -2372 -2016 -2371
rect -2016 -2377 -2009 -2372
rect -2003 -2377 -1997 -2372
rect -1987 -2380 -1983 -2355
rect -1970 -2356 -1952 -2351
rect -1944 -2356 -1884 -2351
rect -1853 -2330 -1841 -2326
rect -1812 -2324 -1785 -2321
rect -1812 -2328 -1809 -2324
rect -1805 -2328 -1792 -2324
rect -1788 -2328 -1785 -2324
rect -1812 -2330 -1785 -2328
rect -1853 -2342 -1849 -2330
rect -1804 -2338 -1800 -2330
rect -1699 -2332 -1672 -2329
rect -1699 -2336 -1696 -2332
rect -1692 -2336 -1679 -2332
rect -1675 -2336 -1672 -2332
rect -1699 -2338 -1672 -2336
rect -1944 -2368 -1940 -2356
rect -1877 -2368 -1868 -2367
rect -1870 -2372 -1868 -2368
rect -1845 -2368 -1841 -2361
rect -1796 -2368 -1792 -2358
rect -1691 -2350 -1687 -2338
rect -1845 -2373 -1804 -2368
rect -1796 -2373 -1703 -2368
rect -1845 -2376 -1841 -2373
rect -1796 -2376 -1792 -2373
rect -1952 -2385 -1948 -2379
rect -1860 -2380 -1823 -2376
rect -1960 -2386 -1933 -2385
rect -1860 -2386 -1856 -2380
rect -1827 -2386 -1823 -2380
rect -1960 -2390 -1959 -2386
rect -1955 -2390 -1938 -2386
rect -1934 -2390 -1933 -2386
rect -1960 -2391 -1933 -2390
rect -1708 -2378 -1691 -2373
rect -1683 -2382 -1679 -2370
rect -1691 -2386 -1679 -2382
rect -1650 -2380 -1623 -2377
rect -1650 -2384 -1647 -2380
rect -1643 -2384 -1630 -2380
rect -1626 -2384 -1623 -2380
rect -1650 -2386 -1623 -2384
rect -1804 -2396 -1800 -2386
rect -1995 -2406 -1991 -2400
rect -1868 -2403 -1864 -2396
rect -1835 -2403 -1831 -2396
rect -1812 -2397 -1785 -2396
rect -1812 -2401 -1811 -2397
rect -1807 -2401 -1790 -2397
rect -1786 -2401 -1785 -2397
rect -1812 -2402 -1785 -2401
rect -1691 -2398 -1687 -2386
rect -1642 -2394 -1638 -2386
rect -1876 -2404 -1849 -2403
rect -2003 -2407 -1976 -2406
rect -2003 -2411 -2002 -2407
rect -1998 -2411 -1981 -2407
rect -1977 -2411 -1976 -2407
rect -1876 -2408 -1875 -2404
rect -1871 -2408 -1854 -2404
rect -1850 -2408 -1849 -2404
rect -1876 -2409 -1849 -2408
rect -1843 -2404 -1816 -2403
rect -1843 -2408 -1842 -2404
rect -1838 -2408 -1821 -2404
rect -1817 -2408 -1816 -2404
rect -1843 -2409 -1816 -2408
rect -2003 -2412 -1976 -2411
rect -1574 -2406 -1569 -2249
rect -1541 -2388 -1514 -2385
rect -1541 -2392 -1538 -2388
rect -1534 -2392 -1521 -2388
rect -1517 -2392 -1514 -2388
rect -1541 -2394 -1514 -2392
rect -1533 -2406 -1529 -2394
rect -1731 -2428 -1706 -2423
rect -1683 -2424 -1679 -2417
rect -1634 -2424 -1630 -2414
rect -1731 -2447 -1726 -2428
rect -1683 -2429 -1642 -2424
rect -1634 -2429 -1553 -2424
rect -1683 -2432 -1679 -2429
rect -1634 -2432 -1630 -2429
rect -1698 -2436 -1661 -2432
rect -1698 -2442 -1694 -2436
rect -1665 -2442 -1661 -2436
rect -2046 -2452 -1726 -2447
rect -1558 -2434 -1533 -2429
rect -1525 -2438 -1521 -2426
rect -1533 -2442 -1521 -2438
rect -1492 -2436 -1465 -2433
rect -1492 -2440 -1489 -2436
rect -1485 -2440 -1472 -2436
rect -1468 -2440 -1465 -2436
rect -1492 -2442 -1465 -2440
rect -1642 -2452 -1638 -2442
rect -1706 -2459 -1702 -2452
rect -1673 -2459 -1669 -2452
rect -1650 -2453 -1623 -2452
rect -1650 -2457 -1649 -2453
rect -1645 -2457 -1628 -2453
rect -1624 -2457 -1623 -2453
rect -1650 -2458 -1623 -2457
rect -1533 -2454 -1529 -2442
rect -1484 -2450 -1480 -2442
rect -1714 -2460 -1687 -2459
rect -1714 -2464 -1713 -2460
rect -1709 -2464 -1692 -2460
rect -1688 -2464 -1687 -2460
rect -1714 -2465 -1687 -2464
rect -1681 -2460 -1654 -2459
rect -1681 -2464 -1680 -2460
rect -1676 -2464 -1659 -2460
rect -1655 -2464 -1654 -2460
rect -1681 -2465 -1654 -2464
rect -1375 -2464 -1348 -2461
rect -1375 -2468 -1372 -2464
rect -1368 -2468 -1355 -2464
rect -1351 -2468 -1348 -2464
rect -1375 -2470 -1348 -2468
rect -1553 -2483 -1548 -2479
rect -1557 -2484 -1548 -2483
rect -1525 -2480 -1521 -2473
rect -1476 -2480 -1472 -2470
rect -1525 -2485 -1484 -2480
rect -1476 -2485 -1385 -2480
rect -1525 -2488 -1521 -2485
rect -1476 -2488 -1472 -2485
rect -1540 -2492 -1503 -2488
rect -1540 -2498 -1536 -2492
rect -1507 -2498 -1503 -2492
rect -1484 -2508 -1480 -2498
rect -1390 -2505 -1385 -2485
rect -1367 -2482 -1363 -2470
rect -1548 -2515 -1544 -2508
rect -1515 -2515 -1511 -2508
rect -1492 -2509 -1465 -2508
rect -1492 -2513 -1491 -2509
rect -1487 -2513 -1470 -2509
rect -1466 -2513 -1465 -2509
rect -1390 -2510 -1367 -2505
rect -1492 -2514 -1465 -2513
rect -1359 -2514 -1355 -2502
rect -1556 -2516 -1529 -2515
rect -1556 -2520 -1555 -2516
rect -1551 -2520 -1534 -2516
rect -1530 -2520 -1529 -2516
rect -1556 -2521 -1529 -2520
rect -1523 -2516 -1496 -2515
rect -1523 -2520 -1522 -2516
rect -1518 -2520 -1501 -2516
rect -1497 -2520 -1496 -2516
rect -1523 -2521 -1496 -2520
rect -1367 -2518 -1355 -2514
rect -1326 -2512 -1299 -2509
rect -1326 -2516 -1323 -2512
rect -1319 -2516 -1306 -2512
rect -1302 -2516 -1299 -2512
rect -1326 -2518 -1299 -2516
rect -1367 -2530 -1363 -2518
rect -1318 -2526 -1314 -2518
rect -1385 -2560 -1382 -2555
rect -1359 -2556 -1355 -2549
rect -1310 -2556 -1306 -2546
rect -1359 -2561 -1318 -2556
rect -1310 -2561 -1297 -2556
rect -1359 -2564 -1355 -2561
rect -1310 -2564 -1306 -2561
rect -1374 -2568 -1337 -2564
rect -1374 -2574 -1370 -2568
rect -1341 -2574 -1337 -2568
rect -1318 -2584 -1314 -2574
rect -1382 -2591 -1378 -2584
rect -1349 -2591 -1345 -2584
rect -1326 -2585 -1299 -2584
rect -1326 -2589 -1325 -2585
rect -1321 -2589 -1304 -2585
rect -1300 -2589 -1299 -2585
rect -1326 -2590 -1299 -2589
rect -1390 -2592 -1363 -2591
rect -1390 -2596 -1389 -2592
rect -1385 -2596 -1368 -2592
rect -1364 -2596 -1363 -2592
rect -1390 -2597 -1363 -2596
rect -1357 -2592 -1330 -2591
rect -1357 -2596 -1356 -2592
rect -1352 -2596 -1335 -2592
rect -1331 -2596 -1330 -2592
rect -1357 -2597 -1330 -2596
rect -2682 -2732 -2381 -2727
rect -2974 -2871 -2658 -2867
rect -3006 -2922 -2972 -2917
rect -2977 -2952 -2972 -2922
rect -2662 -2940 -2658 -2871
rect -2662 -2944 -2657 -2940
rect -2386 -2952 -2381 -2732
rect -2368 -2843 -1605 -2838
rect -2977 -2957 -2328 -2952
rect -3038 -2980 -3011 -2977
rect -3178 -2987 -3143 -2982
rect -3038 -2984 -3035 -2980
rect -3031 -2984 -3018 -2980
rect -3014 -2984 -3011 -2980
rect -3038 -2986 -3011 -2984
rect -3178 -2991 -3172 -2990
rect -3178 -2995 -3177 -2991
rect -3173 -2995 -3172 -2991
rect -3178 -2998 -3172 -2995
rect -3143 -2998 -3138 -2987
rect -3093 -2993 -3084 -2990
rect -3093 -2997 -3091 -2993
rect -3087 -2997 -3084 -2993
rect -3093 -2998 -3084 -2997
rect -3178 -3002 -3166 -2998
rect -3178 -3012 -3172 -3002
rect -3108 -3002 -3084 -2998
rect -3030 -2994 -3026 -2986
rect -3143 -3010 -3128 -3006
rect -3093 -3010 -3084 -3002
rect -3058 -3006 -3045 -3002
rect -3058 -3009 -3054 -3006
rect -3178 -3016 -3177 -3012
rect -3173 -3016 -3172 -3012
rect -3178 -3017 -3172 -3016
rect -3143 -3020 -3138 -3010
rect -3093 -3014 -3091 -3010
rect -3087 -3014 -3084 -3010
rect -3093 -3017 -3084 -3014
rect -3066 -3020 -3062 -3017
rect -3114 -3024 -3062 -3020
rect -3114 -3029 -3110 -3024
rect -3178 -3034 -3110 -3029
rect -3178 -3042 -3172 -3041
rect -3178 -3046 -3177 -3042
rect -3173 -3046 -3172 -3042
rect -3178 -3049 -3172 -3046
rect -3143 -3049 -3138 -3034
rect -3058 -3040 -3054 -3017
rect -3051 -3024 -3045 -3006
rect -3022 -3024 -3018 -3014
rect -2977 -3024 -2972 -2957
rect -2932 -2969 -2878 -2966
rect -2932 -2973 -2929 -2969
rect -2925 -2973 -2912 -2969
rect -2908 -2973 -2902 -2969
rect -2898 -2973 -2885 -2969
rect -2881 -2973 -2878 -2969
rect -2932 -2975 -2878 -2973
rect -2763 -2968 -2709 -2965
rect -2763 -2972 -2760 -2968
rect -2756 -2972 -2743 -2968
rect -2739 -2972 -2733 -2968
rect -2729 -2972 -2716 -2968
rect -2712 -2972 -2709 -2968
rect -2763 -2974 -2709 -2972
rect -2924 -3000 -2920 -2975
rect -2889 -3000 -2885 -2975
rect -3051 -3029 -3030 -3024
rect -3022 -3029 -2972 -3024
rect -3022 -3032 -3018 -3029
rect -3093 -3044 -3084 -3041
rect -3093 -3048 -3091 -3044
rect -3087 -3048 -3084 -3044
rect -3093 -3049 -3084 -3048
rect -3178 -3053 -3166 -3049
rect -3178 -3063 -3172 -3053
rect -3108 -3053 -3084 -3049
rect -3143 -3061 -3128 -3057
rect -3093 -3061 -3084 -3053
rect -3178 -3067 -3177 -3063
rect -3173 -3067 -3172 -3063
rect -3178 -3068 -3172 -3067
rect -3143 -3072 -3138 -3061
rect -3093 -3065 -3091 -3061
rect -3087 -3065 -3084 -3061
rect -3093 -3068 -3084 -3065
rect -3066 -3072 -3062 -3050
rect -3030 -3052 -3026 -3042
rect -3038 -3053 -3011 -3052
rect -3038 -3057 -3037 -3053
rect -3033 -3057 -3016 -3053
rect -3012 -3057 -3011 -3053
rect -3038 -3058 -3011 -3057
rect -3143 -3075 -3062 -3072
rect -3165 -3230 -3111 -3227
rect -3165 -3234 -3162 -3230
rect -3158 -3234 -3145 -3230
rect -3141 -3234 -3135 -3230
rect -3131 -3234 -3118 -3230
rect -3114 -3234 -3111 -3230
rect -3165 -3236 -3111 -3234
rect -3157 -3261 -3153 -3236
rect -3122 -3261 -3118 -3236
rect -3170 -3303 -3157 -3298
rect -3149 -3301 -3145 -3281
rect -3130 -3301 -3126 -3281
rect -3118 -3297 -3111 -3293
rect -3170 -3308 -3165 -3303
rect -3149 -3305 -3126 -3301
rect -3116 -3305 -3111 -3297
rect -3103 -3300 -3076 -3297
rect -3103 -3304 -3100 -3300
rect -3096 -3304 -3083 -3300
rect -3079 -3304 -3076 -3300
rect -3170 -3313 -3139 -3308
rect -3170 -3326 -3165 -3313
rect -3178 -3329 -3165 -3326
rect -3130 -3325 -3126 -3305
rect -3103 -3306 -3076 -3304
rect -3095 -3311 -3091 -3306
rect -3130 -3331 -3107 -3325
rect -3130 -3335 -3126 -3331
rect -3138 -3361 -3134 -3355
rect -3113 -3361 -3107 -3331
rect -2977 -3332 -2972 -3029
rect -2937 -3042 -2924 -3037
rect -2916 -3040 -2912 -3020
rect -2755 -2999 -2751 -2974
rect -2720 -2999 -2716 -2974
rect -2897 -3040 -2893 -3020
rect -2885 -3036 -2878 -3032
rect -2937 -3047 -2932 -3042
rect -2916 -3044 -2893 -3040
rect -2883 -3044 -2878 -3036
rect -2870 -3039 -2843 -3036
rect -2870 -3043 -2867 -3039
rect -2863 -3043 -2850 -3039
rect -2846 -3043 -2843 -3039
rect -2937 -3052 -2906 -3047
rect -2937 -3068 -2932 -3052
rect -2897 -3064 -2893 -3044
rect -2870 -3045 -2843 -3043
rect -2768 -3041 -2755 -3036
rect -2747 -3039 -2743 -3019
rect -2728 -3039 -2724 -3019
rect -2716 -3035 -2709 -3031
rect -2862 -3050 -2858 -3045
rect -2768 -3046 -2763 -3041
rect -2747 -3043 -2724 -3039
rect -2714 -3043 -2709 -3035
rect -2701 -3038 -2674 -3035
rect -2701 -3042 -2698 -3038
rect -2694 -3042 -2681 -3038
rect -2677 -3042 -2674 -3038
rect -2897 -3070 -2874 -3064
rect -2897 -3074 -2893 -3070
rect -2905 -3100 -2901 -3094
rect -2880 -3100 -2874 -3070
rect -2768 -3051 -2737 -3046
rect -2768 -3061 -2763 -3051
rect -2728 -3063 -2724 -3043
rect -2701 -3044 -2674 -3042
rect -2693 -3049 -2689 -3044
rect -2728 -3069 -2705 -3063
rect -2728 -3073 -2724 -3069
rect -2854 -3100 -2850 -3090
rect -2736 -3099 -2732 -3093
rect -2711 -3099 -2705 -3069
rect -2685 -3099 -2681 -3089
rect -2662 -3099 -2657 -2979
rect -2636 -3059 -2631 -2957
rect -2599 -2966 -2545 -2963
rect -2599 -2970 -2596 -2966
rect -2592 -2970 -2579 -2966
rect -2575 -2970 -2569 -2966
rect -2565 -2970 -2552 -2966
rect -2548 -2970 -2545 -2966
rect -2599 -2972 -2545 -2970
rect -2459 -2968 -2405 -2965
rect -2459 -2972 -2456 -2968
rect -2452 -2972 -2439 -2968
rect -2435 -2972 -2429 -2968
rect -2425 -2972 -2412 -2968
rect -2408 -2972 -2405 -2968
rect -2591 -2997 -2587 -2972
rect -2556 -2997 -2552 -2972
rect -2459 -2974 -2405 -2972
rect -2604 -3039 -2591 -3034
rect -2583 -3037 -2579 -3017
rect -2451 -2999 -2447 -2974
rect -2416 -2999 -2412 -2974
rect -2564 -3037 -2560 -3017
rect -2552 -3033 -2545 -3029
rect -2604 -3044 -2599 -3039
rect -2583 -3041 -2560 -3037
rect -2550 -3041 -2545 -3033
rect -2537 -3036 -2510 -3033
rect -2537 -3040 -2534 -3036
rect -2530 -3040 -2517 -3036
rect -2513 -3040 -2510 -3036
rect -2604 -3049 -2573 -3044
rect -2604 -3059 -2599 -3049
rect -2636 -3064 -2599 -3059
rect -2564 -3061 -2560 -3041
rect -2537 -3042 -2510 -3040
rect -2464 -3041 -2451 -3036
rect -2443 -3039 -2439 -3019
rect -2424 -3039 -2420 -3019
rect -2412 -3035 -2405 -3031
rect -2529 -3047 -2525 -3042
rect -2464 -3046 -2459 -3041
rect -2443 -3043 -2420 -3039
rect -2410 -3043 -2405 -3035
rect -2397 -3038 -2370 -3035
rect -2397 -3042 -2394 -3038
rect -2390 -3042 -2377 -3038
rect -2373 -3042 -2370 -3038
rect -2564 -3067 -2541 -3061
rect -2564 -3071 -2560 -3067
rect -2572 -3097 -2568 -3091
rect -2547 -3097 -2541 -3067
rect -2464 -3051 -2433 -3046
rect -2464 -3062 -2459 -3051
rect -2471 -3067 -2459 -3062
rect -2424 -3063 -2420 -3043
rect -2397 -3044 -2370 -3042
rect -2389 -3049 -2385 -3044
rect -2424 -3069 -2401 -3063
rect -2424 -3073 -2420 -3069
rect -2521 -3097 -2517 -3087
rect -2905 -3104 -2893 -3100
rect -2923 -3126 -2919 -3121
rect -2913 -3126 -2907 -3121
rect -2897 -3129 -2893 -3104
rect -2880 -3105 -2862 -3100
rect -2854 -3105 -2757 -3100
rect -2736 -3103 -2724 -3099
rect -2854 -3117 -2850 -3105
rect -2763 -3120 -2757 -3105
rect -2763 -3125 -2750 -3120
rect -2744 -3125 -2738 -3120
rect -2728 -3128 -2724 -3103
rect -2711 -3104 -2693 -3099
rect -2685 -3104 -2593 -3099
rect -2572 -3101 -2560 -3097
rect -2685 -3116 -2681 -3104
rect -2862 -3134 -2858 -3128
rect -2870 -3135 -2843 -3134
rect -2870 -3139 -2869 -3135
rect -2865 -3139 -2848 -3135
rect -2844 -3139 -2843 -3135
rect -2870 -3140 -2843 -3139
rect -2599 -3118 -2593 -3104
rect -2599 -3123 -2586 -3118
rect -2580 -3123 -2574 -3118
rect -2564 -3126 -2560 -3101
rect -2547 -3102 -2529 -3097
rect -2521 -3102 -2481 -3097
rect -2521 -3114 -2517 -3102
rect -2693 -3133 -2689 -3127
rect -2701 -3134 -2674 -3133
rect -2701 -3138 -2700 -3134
rect -2696 -3138 -2679 -3134
rect -2675 -3138 -2674 -3134
rect -2701 -3139 -2674 -3138
rect -2529 -3131 -2525 -3125
rect -2537 -3132 -2510 -3131
rect -2537 -3136 -2536 -3132
rect -2532 -3136 -2515 -3132
rect -2511 -3136 -2510 -3132
rect -2537 -3137 -2510 -3136
rect -2905 -3155 -2901 -3149
rect -2736 -3154 -2732 -3148
rect -2572 -3152 -2568 -3146
rect -2580 -3153 -2553 -3152
rect -2744 -3155 -2717 -3154
rect -2913 -3156 -2886 -3155
rect -2913 -3160 -2912 -3156
rect -2908 -3160 -2891 -3156
rect -2887 -3160 -2886 -3156
rect -2744 -3159 -2743 -3155
rect -2739 -3159 -2722 -3155
rect -2718 -3159 -2717 -3155
rect -2580 -3157 -2579 -3153
rect -2575 -3157 -2558 -3153
rect -2554 -3157 -2553 -3153
rect -2580 -3158 -2553 -3157
rect -2744 -3160 -2717 -3159
rect -2913 -3161 -2886 -3160
rect -2486 -3330 -2481 -3102
rect -2432 -3099 -2428 -3093
rect -2407 -3099 -2401 -3069
rect -2333 -3075 -2328 -2957
rect -2308 -2981 -2254 -2978
rect -2308 -2985 -2305 -2981
rect -2301 -2985 -2288 -2981
rect -2284 -2985 -2278 -2981
rect -2274 -2985 -2261 -2981
rect -2257 -2985 -2254 -2981
rect -2308 -2987 -2254 -2985
rect -2300 -3012 -2296 -2987
rect -2265 -3012 -2261 -2987
rect -2313 -3054 -2300 -3049
rect -2292 -3052 -2288 -3032
rect -1998 -3023 -1971 -3020
rect -1998 -3027 -1995 -3023
rect -1991 -3027 -1978 -3023
rect -1974 -3027 -1971 -3023
rect -1998 -3029 -1971 -3027
rect -2273 -3052 -2269 -3032
rect -1990 -3041 -1986 -3029
rect -2261 -3048 -2254 -3044
rect -2313 -3059 -2308 -3054
rect -2292 -3056 -2269 -3052
rect -2259 -3056 -2254 -3048
rect -2246 -3051 -2219 -3048
rect -2246 -3055 -2243 -3051
rect -2239 -3055 -2226 -3051
rect -2222 -3055 -2219 -3051
rect -2313 -3064 -2282 -3059
rect -2313 -3075 -2308 -3064
rect -2333 -3080 -2308 -3075
rect -2273 -3076 -2269 -3056
rect -2246 -3057 -2219 -3055
rect -2238 -3062 -2234 -3057
rect -2273 -3082 -2250 -3076
rect -2273 -3086 -2269 -3082
rect -2381 -3099 -2377 -3089
rect -2432 -3103 -2420 -3099
rect -2450 -3125 -2446 -3120
rect -2440 -3125 -2434 -3120
rect -2424 -3128 -2420 -3103
rect -2407 -3104 -2389 -3099
rect -2381 -3104 -2350 -3099
rect -2343 -3104 -2302 -3099
rect -2381 -3116 -2377 -3104
rect -2389 -3133 -2385 -3127
rect -2307 -3132 -2302 -3104
rect -2281 -3112 -2277 -3106
rect -2256 -3112 -2250 -3082
rect -2230 -3112 -2226 -3102
rect -2209 -3064 -2011 -3061
rect -2209 -3066 -1990 -3064
rect -2209 -3112 -2204 -3066
rect -2281 -3116 -2269 -3112
rect -2308 -3133 -2302 -3132
rect -2397 -3134 -2370 -3133
rect -2397 -3138 -2396 -3134
rect -2392 -3138 -2375 -3134
rect -2371 -3138 -2370 -3134
rect -2308 -3138 -2295 -3133
rect -2289 -3138 -2283 -3133
rect -2397 -3139 -2370 -3138
rect -2273 -3141 -2269 -3116
rect -2256 -3117 -2238 -3112
rect -2230 -3117 -2204 -3112
rect -2230 -3129 -2226 -3117
rect -2432 -3154 -2428 -3148
rect -2440 -3155 -2413 -3154
rect -2440 -3159 -2439 -3155
rect -2435 -3159 -2418 -3155
rect -2414 -3159 -2413 -3155
rect -2440 -3160 -2413 -3159
rect -2238 -3146 -2234 -3140
rect -2246 -3147 -2219 -3146
rect -2246 -3151 -2245 -3147
rect -2241 -3151 -2224 -3147
rect -2220 -3151 -2219 -3147
rect -2246 -3152 -2219 -3151
rect -2281 -3167 -2277 -3161
rect -2289 -3168 -2262 -3167
rect -2289 -3172 -2288 -3168
rect -2284 -3172 -2267 -3168
rect -2263 -3172 -2262 -3168
rect -2289 -3173 -2262 -3172
rect -2184 -3280 -2179 -3066
rect -2016 -3069 -1990 -3066
rect -1982 -3073 -1978 -3061
rect -1990 -3077 -1978 -3073
rect -1949 -3071 -1922 -3068
rect -1949 -3075 -1946 -3071
rect -1942 -3075 -1929 -3071
rect -1925 -3075 -1922 -3071
rect -1949 -3077 -1922 -3075
rect -1990 -3089 -1986 -3077
rect -1941 -3085 -1937 -3077
rect -2010 -3119 -2005 -3114
rect -1982 -3115 -1978 -3108
rect -1933 -3115 -1929 -3105
rect -1982 -3120 -1941 -3115
rect -1933 -3120 -1910 -3115
rect -1982 -3123 -1978 -3120
rect -1933 -3123 -1929 -3120
rect -1997 -3127 -1960 -3123
rect -1997 -3133 -1993 -3127
rect -1964 -3133 -1960 -3127
rect -1941 -3143 -1937 -3133
rect -2005 -3150 -2001 -3143
rect -1972 -3150 -1968 -3143
rect -1949 -3144 -1922 -3143
rect -1949 -3148 -1948 -3144
rect -1944 -3148 -1927 -3144
rect -1923 -3148 -1922 -3144
rect -1949 -3149 -1922 -3148
rect -2013 -3151 -1986 -3150
rect -2013 -3155 -2012 -3151
rect -2008 -3155 -1991 -3151
rect -1987 -3155 -1986 -3151
rect -2013 -3156 -1986 -3155
rect -1980 -3151 -1953 -3150
rect -1980 -3155 -1979 -3151
rect -1975 -3155 -1958 -3151
rect -1954 -3155 -1953 -3151
rect -1980 -3156 -1953 -3155
rect -2145 -3185 -2091 -3182
rect -2145 -3189 -2142 -3185
rect -2138 -3189 -2125 -3185
rect -2121 -3189 -2115 -3185
rect -2111 -3189 -2098 -3185
rect -2094 -3189 -2091 -3185
rect -2145 -3191 -2091 -3189
rect -2137 -3216 -2133 -3191
rect -2102 -3216 -2098 -3191
rect -2150 -3258 -2137 -3253
rect -2129 -3256 -2125 -3236
rect -2110 -3256 -2106 -3236
rect -2098 -3252 -2091 -3248
rect -2150 -3263 -2145 -3258
rect -2129 -3260 -2106 -3256
rect -2096 -3260 -2091 -3252
rect -2083 -3255 -2056 -3252
rect -2083 -3259 -2080 -3255
rect -2076 -3259 -2063 -3255
rect -2059 -3259 -2056 -3255
rect -2150 -3268 -2119 -3263
rect -2150 -3280 -2145 -3268
rect -2184 -3285 -2145 -3280
rect -2110 -3280 -2106 -3260
rect -2083 -3261 -2056 -3259
rect -2075 -3266 -2071 -3261
rect -2110 -3286 -2087 -3280
rect -2110 -3290 -2106 -3286
rect -2118 -3316 -2114 -3310
rect -2093 -3316 -2087 -3286
rect -1915 -3273 -1910 -3120
rect -1864 -3233 -1837 -3230
rect -1864 -3237 -1861 -3233
rect -1857 -3237 -1844 -3233
rect -1840 -3237 -1837 -3233
rect -1864 -3239 -1837 -3237
rect -1856 -3251 -1852 -3239
rect -1915 -3274 -1868 -3273
rect -1915 -3278 -1856 -3274
rect -1873 -3279 -1856 -3278
rect -1848 -3283 -1844 -3271
rect -2067 -3316 -2063 -3306
rect -1856 -3287 -1844 -3283
rect -1815 -3281 -1788 -3278
rect -1815 -3285 -1812 -3281
rect -1808 -3285 -1795 -3281
rect -1791 -3285 -1788 -3281
rect -1815 -3287 -1788 -3285
rect -1856 -3299 -1852 -3287
rect -1807 -3295 -1803 -3287
rect -2118 -3320 -2106 -3316
rect -2977 -3337 -2543 -3332
rect -2486 -3335 -2168 -3330
rect -2163 -3335 -2139 -3330
rect -2148 -3337 -2139 -3335
rect -2148 -3342 -2132 -3337
rect -2126 -3342 -2120 -3337
rect -2148 -3343 -2139 -3342
rect -2110 -3345 -2106 -3320
rect -2093 -3321 -2075 -3316
rect -2067 -3321 -1903 -3316
rect -2067 -3333 -2063 -3321
rect -1908 -3323 -1903 -3321
rect -1908 -3324 -1877 -3323
rect -1908 -3328 -1871 -3324
rect -1880 -3329 -1871 -3328
rect -1848 -3325 -1844 -3318
rect -1799 -3325 -1795 -3315
rect -1848 -3330 -1807 -3325
rect -1799 -3330 -1749 -3325
rect -1848 -3333 -1844 -3330
rect -1799 -3333 -1795 -3330
rect -3087 -3361 -3083 -3351
rect -3138 -3365 -3126 -3361
rect -3165 -3382 -3159 -3365
rect -3165 -3387 -3152 -3382
rect -3146 -3387 -3140 -3382
rect -3130 -3390 -3126 -3365
rect -3113 -3366 -3095 -3361
rect -3087 -3366 -2156 -3361
rect -3087 -3378 -3083 -3366
rect -3095 -3395 -3091 -3389
rect -3103 -3396 -3076 -3395
rect -3103 -3400 -3102 -3396
rect -3098 -3400 -3081 -3396
rect -3077 -3400 -3076 -3396
rect -3103 -3401 -3076 -3400
rect -2161 -3396 -2156 -3366
rect -1863 -3337 -1826 -3333
rect -1863 -3343 -1859 -3337
rect -1830 -3343 -1826 -3337
rect -2075 -3350 -2071 -3344
rect -2083 -3351 -2056 -3350
rect -2083 -3355 -2082 -3351
rect -2078 -3355 -2061 -3351
rect -2057 -3355 -2056 -3351
rect -2083 -3356 -2056 -3355
rect -1807 -3353 -1803 -3343
rect -1871 -3360 -1867 -3353
rect -1838 -3360 -1834 -3353
rect -1815 -3354 -1788 -3353
rect -1815 -3358 -1814 -3354
rect -1810 -3358 -1793 -3354
rect -1789 -3358 -1788 -3354
rect -1815 -3359 -1788 -3358
rect -1879 -3361 -1852 -3360
rect -1879 -3365 -1878 -3361
rect -1874 -3365 -1857 -3361
rect -1853 -3365 -1852 -3361
rect -2118 -3371 -2114 -3365
rect -1879 -3366 -1852 -3365
rect -1846 -3361 -1819 -3360
rect -1846 -3365 -1845 -3361
rect -1841 -3365 -1824 -3361
rect -1820 -3365 -1819 -3361
rect -1846 -3366 -1819 -3365
rect -2126 -3372 -2099 -3371
rect -2126 -3376 -2125 -3372
rect -2121 -3376 -2104 -3372
rect -2100 -3376 -2099 -3372
rect -2126 -3377 -2099 -3376
rect -2161 -3401 -1803 -3396
rect -3138 -3416 -3134 -3410
rect -3146 -3417 -3119 -3416
rect -3146 -3421 -3145 -3417
rect -3141 -3421 -3124 -3417
rect -3120 -3421 -3119 -3417
rect -3146 -3422 -3119 -3421
rect -1808 -3484 -1803 -3401
rect -1754 -3434 -1749 -3330
rect -1717 -3393 -1690 -3390
rect -1717 -3397 -1714 -3393
rect -1710 -3397 -1697 -3393
rect -1693 -3397 -1690 -3393
rect -1717 -3399 -1690 -3397
rect -1709 -3411 -1705 -3399
rect -1754 -3439 -1709 -3434
rect -1701 -3443 -1697 -3431
rect -1709 -3447 -1697 -3443
rect -1668 -3441 -1641 -3438
rect -1668 -3445 -1665 -3441
rect -1661 -3445 -1648 -3441
rect -1644 -3445 -1641 -3441
rect -1668 -3447 -1641 -3445
rect -1610 -3445 -1605 -2843
rect -1499 -3424 -1495 -3414
rect -1559 -3437 -1518 -3432
rect -1559 -3445 -1554 -3437
rect -1709 -3459 -1705 -3447
rect -1660 -3455 -1656 -3447
rect -1610 -3450 -1554 -3445
rect -1523 -3451 -1518 -3437
rect -1523 -3452 -1507 -3451
rect -1523 -3456 -1498 -3452
rect -1808 -3489 -1752 -3484
rect -1745 -3489 -1724 -3484
rect -1701 -3485 -1697 -3478
rect -1652 -3485 -1648 -3475
rect -1509 -3466 -1506 -3456
rect -1491 -3457 -1487 -3444
rect -1509 -3479 -1506 -3471
rect -1499 -3472 -1495 -3467
rect -1481 -3472 -1480 -3468
rect -1509 -3483 -1499 -3479
rect -1701 -3490 -1660 -3485
rect -1652 -3490 -1521 -3485
rect -1701 -3493 -1697 -3490
rect -1652 -3493 -1648 -3490
rect -1716 -3497 -1679 -3493
rect -1716 -3503 -1712 -3497
rect -1683 -3503 -1679 -3497
rect -1660 -3513 -1656 -3503
rect -1526 -3508 -1521 -3490
rect -1491 -3506 -1487 -3499
rect -1481 -3506 -1477 -3499
rect -1506 -3508 -1498 -3506
rect -1526 -3510 -1498 -3508
rect -1491 -3510 -1477 -3506
rect -1526 -3513 -1503 -3510
rect -1724 -3520 -1720 -3513
rect -1691 -3520 -1687 -3513
rect -1668 -3514 -1641 -3513
rect -1668 -3518 -1667 -3514
rect -1663 -3518 -1646 -3514
rect -1642 -3518 -1641 -3514
rect -1668 -3519 -1641 -3518
rect -1732 -3521 -1705 -3520
rect -1732 -3525 -1731 -3521
rect -1727 -3525 -1710 -3521
rect -1706 -3525 -1705 -3521
rect -1732 -3526 -1705 -3525
rect -1699 -3521 -1672 -3520
rect -1699 -3525 -1698 -3521
rect -1694 -3525 -1677 -3521
rect -1673 -3525 -1672 -3521
rect -1699 -3526 -1672 -3525
rect -1506 -3530 -1503 -3513
rect -1491 -3511 -1487 -3510
rect -1481 -3511 -1477 -3510
rect -1473 -3506 -1469 -3499
rect -1473 -3510 -1457 -3506
rect -1473 -3511 -1469 -3510
rect -1499 -3522 -1495 -3521
rect -1482 -3526 -1474 -3522
rect -1470 -3526 -1468 -3522
rect -1460 -3530 -1457 -3510
rect -1506 -3533 -1457 -3530
rect -2911 -3742 -2857 -3739
rect -3038 -3748 -3011 -3745
rect -2911 -3746 -2908 -3742
rect -2904 -3746 -2891 -3742
rect -2887 -3746 -2881 -3742
rect -2877 -3746 -2864 -3742
rect -2860 -3746 -2857 -3742
rect -2911 -3748 -2857 -3746
rect -3178 -3755 -3143 -3750
rect -3038 -3752 -3035 -3748
rect -3031 -3752 -3018 -3748
rect -3014 -3752 -3011 -3748
rect -3038 -3754 -3011 -3752
rect -3178 -3759 -3172 -3758
rect -3178 -3763 -3177 -3759
rect -3173 -3763 -3172 -3759
rect -3178 -3766 -3172 -3763
rect -3143 -3766 -3138 -3755
rect -3093 -3761 -3084 -3758
rect -3093 -3765 -3091 -3761
rect -3087 -3765 -3084 -3761
rect -3093 -3766 -3084 -3765
rect -3178 -3770 -3166 -3766
rect -3178 -3780 -3172 -3770
rect -3108 -3770 -3084 -3766
rect -3030 -3762 -3026 -3754
rect -3143 -3778 -3128 -3774
rect -3093 -3778 -3084 -3770
rect -3058 -3774 -3045 -3770
rect -3058 -3777 -3054 -3774
rect -3178 -3784 -3177 -3780
rect -3173 -3784 -3172 -3780
rect -3178 -3785 -3172 -3784
rect -3143 -3788 -3138 -3778
rect -3093 -3782 -3091 -3778
rect -3087 -3782 -3084 -3778
rect -3093 -3785 -3084 -3782
rect -3066 -3788 -3062 -3785
rect -3114 -3792 -3062 -3788
rect -3114 -3797 -3110 -3792
rect -3178 -3802 -3110 -3797
rect -3178 -3810 -3172 -3809
rect -3178 -3814 -3177 -3810
rect -3173 -3814 -3172 -3810
rect -3178 -3817 -3172 -3814
rect -3143 -3817 -3138 -3802
rect -3058 -3808 -3054 -3785
rect -3051 -3792 -3045 -3774
rect -3022 -3792 -3018 -3782
rect -2903 -3773 -2899 -3748
rect -2868 -3773 -2864 -3748
rect -3051 -3797 -3030 -3792
rect -3022 -3797 -2960 -3792
rect -3022 -3800 -3018 -3797
rect -3093 -3812 -3084 -3809
rect -3093 -3816 -3091 -3812
rect -3087 -3816 -3084 -3812
rect -3093 -3817 -3084 -3816
rect -3178 -3821 -3166 -3817
rect -3178 -3831 -3172 -3821
rect -3108 -3821 -3084 -3817
rect -3143 -3829 -3128 -3825
rect -3093 -3829 -3084 -3821
rect -3178 -3835 -3177 -3831
rect -3173 -3835 -3172 -3831
rect -3178 -3836 -3172 -3835
rect -3143 -3840 -3138 -3829
rect -3093 -3833 -3091 -3829
rect -3087 -3833 -3084 -3829
rect -3093 -3836 -3084 -3833
rect -3066 -3840 -3062 -3818
rect -3030 -3820 -3026 -3810
rect -3038 -3821 -3011 -3820
rect -3038 -3825 -3037 -3821
rect -3033 -3825 -3016 -3821
rect -3012 -3825 -3011 -3821
rect -3038 -3826 -3011 -3825
rect -3143 -3843 -3062 -3840
rect -3171 -4079 -3117 -4076
rect -3171 -4083 -3168 -4079
rect -3164 -4083 -3151 -4079
rect -3147 -4083 -3141 -4079
rect -3137 -4083 -3124 -4079
rect -3120 -4083 -3117 -4079
rect -3171 -4085 -3117 -4083
rect -3163 -4110 -3159 -4085
rect -3128 -4110 -3124 -4085
rect -3176 -4152 -3163 -4147
rect -3155 -4150 -3151 -4130
rect -3136 -4150 -3132 -4130
rect -3124 -4146 -3117 -4142
rect -3176 -4157 -3171 -4152
rect -3155 -4154 -3132 -4150
rect -3122 -4154 -3117 -4146
rect -3109 -4149 -3082 -4146
rect -3109 -4153 -3106 -4149
rect -3102 -4153 -3089 -4149
rect -3085 -4153 -3082 -4149
rect -3176 -4162 -3145 -4157
rect -3176 -4175 -3171 -4162
rect -3184 -4178 -3171 -4175
rect -3136 -4174 -3132 -4154
rect -3109 -4155 -3082 -4153
rect -3101 -4160 -3097 -4155
rect -3136 -4180 -3113 -4174
rect -3136 -4184 -3132 -4180
rect -3144 -4210 -3140 -4204
rect -3119 -4210 -3113 -4180
rect -2992 -4192 -2987 -3797
rect -2965 -3837 -2960 -3797
rect -2916 -3815 -2903 -3810
rect -2895 -3813 -2891 -3793
rect -2876 -3813 -2872 -3793
rect -2864 -3809 -2857 -3805
rect -2916 -3820 -2911 -3815
rect -2895 -3817 -2872 -3813
rect -2862 -3817 -2857 -3809
rect -2849 -3812 -2822 -3809
rect -2849 -3816 -2846 -3812
rect -2842 -3816 -2829 -3812
rect -2825 -3816 -2822 -3812
rect -2916 -3825 -2885 -3820
rect -2916 -3837 -2911 -3825
rect -2965 -3842 -2939 -3837
rect -2934 -3842 -2930 -3837
rect -2925 -3842 -2911 -3837
rect -2876 -3837 -2872 -3817
rect -2849 -3818 -2822 -3816
rect -2841 -3823 -2837 -3818
rect -2876 -3843 -2853 -3837
rect -2876 -3847 -2872 -3843
rect -2884 -3873 -2880 -3867
rect -2859 -3873 -2853 -3843
rect -2833 -3873 -2829 -3863
rect -2953 -3883 -2905 -3876
rect -2884 -3877 -2872 -3873
rect -2912 -3894 -2905 -3883
rect -2912 -3899 -2898 -3894
rect -2892 -3899 -2886 -3894
rect -2876 -3902 -2872 -3877
rect -2859 -3878 -2841 -3873
rect -2833 -3878 -2766 -3873
rect -2833 -3890 -2829 -3878
rect -2841 -3907 -2837 -3901
rect -2849 -3908 -2822 -3907
rect -2849 -3912 -2848 -3908
rect -2844 -3912 -2827 -3908
rect -2823 -3912 -2822 -3908
rect -2849 -3913 -2822 -3912
rect -2884 -3928 -2880 -3922
rect -2771 -3924 -2766 -3878
rect -2745 -3883 -2718 -3880
rect -2745 -3887 -2742 -3883
rect -2738 -3887 -2725 -3883
rect -2721 -3887 -2718 -3883
rect -2745 -3889 -2718 -3887
rect -2737 -3901 -2733 -3889
rect -2892 -3929 -2865 -3928
rect -2771 -3929 -2737 -3924
rect -2892 -3933 -2891 -3929
rect -2887 -3933 -2870 -3929
rect -2866 -3933 -2865 -3929
rect -2729 -3933 -2725 -3921
rect -2892 -3934 -2865 -3933
rect -2737 -3937 -2725 -3933
rect -2696 -3931 -2669 -3928
rect -2696 -3935 -2693 -3931
rect -2689 -3935 -2676 -3931
rect -2672 -3935 -2669 -3931
rect -2696 -3937 -2669 -3935
rect -2910 -3947 -2856 -3944
rect -2910 -3951 -2907 -3947
rect -2903 -3951 -2890 -3947
rect -2886 -3951 -2880 -3947
rect -2876 -3951 -2863 -3947
rect -2859 -3951 -2856 -3947
rect -2910 -3953 -2856 -3951
rect -2737 -3949 -2733 -3937
rect -2688 -3945 -2684 -3937
rect -2902 -3978 -2898 -3953
rect -2867 -3978 -2863 -3953
rect -2915 -4020 -2902 -4015
rect -2894 -4018 -2890 -3998
rect -2789 -3973 -2761 -3972
rect -2789 -3974 -2760 -3973
rect -2789 -3977 -2752 -3974
rect -2875 -4018 -2871 -3998
rect -2863 -4014 -2856 -4010
rect -2915 -4025 -2910 -4020
rect -2894 -4022 -2871 -4018
rect -2861 -4022 -2856 -4014
rect -2848 -4017 -2821 -4014
rect -2848 -4021 -2845 -4017
rect -2841 -4021 -2828 -4017
rect -2824 -4021 -2821 -4017
rect -2915 -4030 -2884 -4025
rect -2915 -4041 -2910 -4030
rect -2918 -4046 -2910 -4041
rect -2875 -4042 -2871 -4022
rect -2848 -4023 -2821 -4021
rect -2840 -4028 -2836 -4023
rect -2875 -4048 -2852 -4042
rect -2875 -4052 -2871 -4048
rect -2883 -4078 -2879 -4072
rect -2858 -4078 -2852 -4048
rect -2832 -4078 -2828 -4068
rect -2789 -4078 -2784 -3977
rect -2766 -3979 -2752 -3977
rect -2729 -3975 -2725 -3968
rect -2680 -3975 -2676 -3965
rect -2729 -3980 -2688 -3975
rect -2680 -3980 -2640 -3975
rect -2729 -3983 -2725 -3980
rect -2680 -3983 -2676 -3980
rect -2744 -3987 -2707 -3983
rect -2744 -3993 -2740 -3987
rect -2711 -3993 -2707 -3987
rect -2688 -4003 -2684 -3993
rect -2752 -4010 -2748 -4003
rect -2719 -4010 -2715 -4003
rect -2696 -4004 -2669 -4003
rect -2696 -4008 -2695 -4004
rect -2691 -4008 -2674 -4004
rect -2670 -4008 -2669 -4004
rect -2696 -4009 -2669 -4008
rect -2760 -4011 -2733 -4010
rect -2760 -4015 -2759 -4011
rect -2755 -4015 -2738 -4011
rect -2734 -4015 -2733 -4011
rect -2760 -4016 -2733 -4015
rect -2727 -4011 -2700 -4010
rect -2727 -4015 -2726 -4011
rect -2722 -4015 -2705 -4011
rect -2701 -4015 -2700 -4011
rect -2727 -4016 -2700 -4015
rect -2645 -4037 -2640 -3980
rect -2599 -3996 -2572 -3993
rect -2599 -4000 -2596 -3996
rect -2592 -4000 -2579 -3996
rect -2575 -4000 -2572 -3996
rect -2599 -4002 -2572 -4000
rect -2591 -4014 -2587 -4002
rect -2645 -4042 -2591 -4037
rect -2583 -4046 -2579 -4034
rect -2417 -4035 -2413 -4025
rect -2883 -4082 -2871 -4078
rect -2904 -4104 -2897 -4099
rect -2891 -4104 -2885 -4099
rect -2875 -4107 -2871 -4082
rect -2858 -4083 -2840 -4078
rect -2832 -4083 -2784 -4078
rect -2591 -4050 -2579 -4046
rect -2550 -4044 -2523 -4041
rect -2550 -4048 -2547 -4044
rect -2543 -4048 -2530 -4044
rect -2526 -4048 -2523 -4044
rect -2550 -4050 -2523 -4048
rect -2591 -4062 -2587 -4050
rect -2542 -4058 -2538 -4050
rect -2832 -4095 -2828 -4083
rect -2615 -4088 -2606 -4087
rect -2659 -4093 -2633 -4088
rect -2623 -4092 -2606 -4088
rect -2583 -4088 -2579 -4081
rect -2534 -4088 -2530 -4078
rect -2422 -4067 -2416 -4063
rect -2409 -4068 -2405 -4055
rect -2427 -4077 -2424 -4068
rect -2623 -4093 -2612 -4092
rect -2583 -4093 -2542 -4088
rect -2534 -4093 -2446 -4088
rect -2840 -4112 -2836 -4106
rect -2848 -4113 -2821 -4112
rect -2848 -4117 -2847 -4113
rect -2843 -4117 -2826 -4113
rect -2822 -4117 -2821 -4113
rect -2848 -4118 -2821 -4117
rect -2883 -4133 -2879 -4127
rect -2891 -4134 -2864 -4133
rect -2891 -4138 -2890 -4134
rect -2886 -4138 -2869 -4134
rect -2865 -4138 -2864 -4134
rect -2891 -4139 -2864 -4138
rect -3093 -4210 -3089 -4200
rect -2659 -4210 -2654 -4093
rect -2583 -4096 -2579 -4093
rect -2534 -4096 -2530 -4093
rect -2598 -4100 -2561 -4096
rect -2598 -4106 -2594 -4100
rect -2565 -4106 -2561 -4100
rect -2542 -4116 -2538 -4106
rect -2606 -4123 -2602 -4116
rect -2573 -4123 -2569 -4116
rect -2550 -4117 -2523 -4116
rect -2550 -4121 -2549 -4117
rect -2545 -4121 -2528 -4117
rect -2524 -4121 -2523 -4117
rect -2550 -4122 -2523 -4121
rect -2451 -4119 -2446 -4093
rect -2427 -4090 -2424 -4082
rect -2417 -4083 -2413 -4078
rect -2399 -4083 -2398 -4079
rect -2427 -4094 -2417 -4090
rect -2409 -4117 -2405 -4110
rect -2399 -4117 -2395 -4110
rect -2424 -4119 -2416 -4117
rect -2451 -4121 -2416 -4119
rect -2409 -4121 -2395 -4117
rect -2614 -4124 -2587 -4123
rect -2614 -4128 -2613 -4124
rect -2609 -4128 -2592 -4124
rect -2588 -4128 -2587 -4124
rect -2614 -4129 -2587 -4128
rect -2581 -4124 -2554 -4123
rect -2451 -4124 -2421 -4121
rect -2581 -4128 -2580 -4124
rect -2576 -4128 -2559 -4124
rect -2555 -4128 -2554 -4124
rect -2581 -4129 -2554 -4128
rect -2424 -4141 -2421 -4124
rect -2409 -4122 -2405 -4121
rect -2399 -4122 -2395 -4121
rect -2391 -4117 -2387 -4110
rect -2391 -4121 -2375 -4117
rect -2391 -4122 -2387 -4121
rect -2417 -4133 -2413 -4132
rect -2400 -4137 -2392 -4133
rect -2388 -4137 -2386 -4133
rect -2378 -4141 -2375 -4121
rect 708 -4135 712 -4125
rect -2424 -4144 -2375 -4141
rect 698 -4167 709 -4163
rect 698 -4177 701 -4167
rect 716 -4168 720 -4155
rect 698 -4190 701 -4182
rect 708 -4183 712 -4178
rect 726 -4183 727 -4179
rect 698 -4194 708 -4190
rect -3144 -4214 -3132 -4210
rect -3171 -4231 -3165 -4214
rect -3171 -4236 -3158 -4231
rect -3152 -4236 -3146 -4231
rect -3136 -4239 -3132 -4214
rect -3119 -4215 -3101 -4210
rect -3093 -4215 -2654 -4210
rect -3093 -4227 -3089 -4215
rect 716 -4217 720 -4210
rect 726 -4217 730 -4210
rect 701 -4221 709 -4217
rect 716 -4221 730 -4217
rect -2992 -4235 -2987 -4231
rect -3101 -4244 -3097 -4238
rect -3109 -4245 -3082 -4244
rect -3109 -4249 -3108 -4245
rect -3104 -4249 -3087 -4245
rect -3083 -4249 -3082 -4245
rect -3109 -4250 -3082 -4249
rect -3144 -4265 -3140 -4259
rect -3152 -4266 -3125 -4265
rect -3152 -4270 -3151 -4266
rect -3147 -4270 -3130 -4266
rect -3126 -4270 -3125 -4266
rect -3152 -4271 -3125 -4270
rect -2991 -4285 -2987 -4235
rect 701 -4241 704 -4221
rect 716 -4222 720 -4221
rect 726 -4222 730 -4221
rect 734 -4217 738 -4210
rect 734 -4221 750 -4217
rect 734 -4222 738 -4221
rect 708 -4233 712 -4232
rect 725 -4237 733 -4233
rect 737 -4237 739 -4233
rect 747 -4241 750 -4221
rect 701 -4244 750 -4241
rect -2991 -4289 -2729 -4285
rect -2954 -4380 -2886 -4373
rect -3060 -4510 -3033 -4507
rect -3200 -4517 -3165 -4512
rect -3060 -4514 -3057 -4510
rect -3053 -4514 -3040 -4510
rect -3036 -4514 -3033 -4510
rect -3060 -4516 -3033 -4514
rect -3200 -4521 -3194 -4520
rect -3200 -4525 -3199 -4521
rect -3195 -4525 -3194 -4521
rect -3200 -4528 -3194 -4525
rect -3165 -4528 -3160 -4517
rect -3115 -4523 -3106 -4520
rect -3115 -4527 -3113 -4523
rect -3109 -4527 -3106 -4523
rect -3115 -4528 -3106 -4527
rect -3200 -4532 -3188 -4528
rect -3200 -4542 -3194 -4532
rect -3130 -4532 -3106 -4528
rect -3052 -4524 -3048 -4516
rect -2999 -4522 -2945 -4519
rect -3165 -4540 -3150 -4536
rect -3115 -4540 -3106 -4532
rect -3080 -4536 -3067 -4532
rect -3080 -4539 -3076 -4536
rect -3200 -4546 -3199 -4542
rect -3195 -4546 -3194 -4542
rect -3200 -4547 -3194 -4546
rect -3165 -4550 -3160 -4540
rect -3115 -4544 -3113 -4540
rect -3109 -4544 -3106 -4540
rect -3115 -4547 -3106 -4544
rect -3088 -4550 -3084 -4547
rect -3136 -4554 -3084 -4550
rect -3136 -4559 -3132 -4554
rect -3200 -4564 -3132 -4559
rect -3200 -4572 -3194 -4571
rect -3200 -4576 -3199 -4572
rect -3195 -4576 -3194 -4572
rect -3200 -4579 -3194 -4576
rect -3165 -4579 -3160 -4564
rect -3080 -4570 -3076 -4547
rect -3073 -4554 -3067 -4536
rect -2999 -4526 -2996 -4522
rect -2992 -4526 -2979 -4522
rect -2975 -4526 -2969 -4522
rect -2965 -4526 -2952 -4522
rect -2948 -4526 -2945 -4522
rect -2999 -4528 -2945 -4526
rect -3044 -4554 -3040 -4544
rect -2991 -4553 -2987 -4528
rect -2956 -4553 -2952 -4528
rect -3073 -4559 -3052 -4554
rect -3044 -4559 -3026 -4554
rect -3044 -4562 -3040 -4559
rect -3115 -4574 -3106 -4571
rect -3115 -4578 -3113 -4574
rect -3109 -4578 -3106 -4574
rect -3115 -4579 -3106 -4578
rect -3200 -4583 -3188 -4579
rect -3200 -4593 -3194 -4583
rect -3130 -4583 -3106 -4579
rect -3165 -4591 -3150 -4587
rect -3115 -4591 -3106 -4583
rect -3200 -4597 -3199 -4593
rect -3195 -4597 -3194 -4593
rect -3200 -4598 -3194 -4597
rect -3165 -4602 -3160 -4591
rect -3115 -4595 -3113 -4591
rect -3109 -4595 -3106 -4591
rect -3115 -4598 -3106 -4595
rect -3088 -4602 -3084 -4580
rect -3052 -4582 -3048 -4572
rect -3031 -4579 -3026 -4559
rect -3060 -4583 -3033 -4582
rect -3060 -4587 -3059 -4583
rect -3055 -4587 -3038 -4583
rect -3034 -4587 -3033 -4583
rect -3060 -4588 -3033 -4587
rect -3030 -4596 -3026 -4579
rect -3165 -4605 -3084 -4602
rect -3031 -4616 -3026 -4596
rect -3004 -4595 -2991 -4590
rect -2983 -4593 -2979 -4573
rect -2964 -4593 -2960 -4573
rect -2952 -4589 -2945 -4585
rect -3004 -4600 -2999 -4595
rect -2983 -4597 -2960 -4593
rect -2950 -4597 -2945 -4589
rect -2937 -4592 -2910 -4589
rect -2937 -4596 -2934 -4592
rect -2930 -4596 -2917 -4592
rect -2913 -4596 -2910 -4592
rect -3004 -4605 -2973 -4600
rect -3004 -4616 -2999 -4605
rect -3031 -4621 -3008 -4616
rect -3003 -4621 -2999 -4616
rect -2964 -4617 -2960 -4597
rect -2937 -4598 -2910 -4596
rect -2929 -4603 -2925 -4598
rect -3168 -4702 -3114 -4699
rect -3168 -4706 -3165 -4702
rect -3161 -4706 -3148 -4702
rect -3144 -4706 -3138 -4702
rect -3134 -4706 -3121 -4702
rect -3117 -4706 -3114 -4702
rect -3168 -4708 -3114 -4706
rect -3160 -4733 -3156 -4708
rect -3125 -4733 -3121 -4708
rect -3173 -4775 -3160 -4770
rect -3152 -4773 -3148 -4753
rect -3133 -4773 -3129 -4753
rect -3121 -4769 -3114 -4765
rect -3173 -4780 -3168 -4775
rect -3152 -4777 -3129 -4773
rect -3119 -4777 -3114 -4769
rect -3106 -4772 -3079 -4769
rect -3106 -4776 -3103 -4772
rect -3099 -4776 -3086 -4772
rect -3082 -4776 -3079 -4772
rect -3173 -4785 -3142 -4780
rect -3173 -4798 -3168 -4785
rect -3181 -4801 -3168 -4798
rect -3133 -4797 -3129 -4777
rect -3106 -4778 -3079 -4776
rect -3098 -4783 -3094 -4778
rect -3133 -4803 -3110 -4797
rect -3133 -4807 -3129 -4803
rect -3141 -4833 -3137 -4827
rect -3116 -4833 -3110 -4803
rect -3031 -4816 -3026 -4621
rect -2964 -4623 -2941 -4617
rect -2964 -4627 -2960 -4623
rect -2972 -4653 -2968 -4647
rect -2947 -4653 -2941 -4623
rect -2921 -4653 -2917 -4643
rect -2972 -4657 -2960 -4653
rect -2999 -4679 -2986 -4674
rect -2980 -4679 -2974 -4674
rect -2999 -4812 -2994 -4679
rect -2964 -4682 -2960 -4657
rect -2947 -4658 -2929 -4653
rect -2921 -4658 -2890 -4653
rect -2921 -4670 -2917 -4658
rect -2929 -4687 -2925 -4681
rect -2937 -4688 -2910 -4687
rect -2937 -4692 -2936 -4688
rect -2932 -4692 -2915 -4688
rect -2911 -4692 -2910 -4688
rect -2937 -4693 -2910 -4692
rect -2972 -4708 -2968 -4702
rect -2980 -4709 -2953 -4708
rect -2980 -4713 -2979 -4709
rect -2975 -4713 -2958 -4709
rect -2954 -4713 -2953 -4709
rect -2980 -4714 -2953 -4713
rect -2895 -4765 -2890 -4658
rect -2851 -4726 -2824 -4723
rect -2851 -4730 -2848 -4726
rect -2844 -4730 -2831 -4726
rect -2827 -4730 -2824 -4726
rect -2851 -4732 -2824 -4730
rect -2843 -4744 -2839 -4732
rect -2895 -4770 -2885 -4765
rect -2878 -4767 -2855 -4765
rect -2878 -4770 -2843 -4767
rect -2860 -4772 -2843 -4770
rect -2835 -4776 -2831 -4764
rect -2733 -4764 -2729 -4289
rect -2609 -4759 -2605 -4751
rect -2733 -4768 -2668 -4764
rect -2843 -4780 -2831 -4776
rect -2802 -4774 -2775 -4771
rect -2802 -4778 -2799 -4774
rect -2795 -4778 -2782 -4774
rect -2778 -4778 -2775 -4774
rect -2802 -4780 -2775 -4778
rect -2843 -4792 -2839 -4780
rect -2794 -4788 -2790 -4780
rect -2672 -4784 -2668 -4768
rect -2672 -4787 -2616 -4784
rect -2672 -4788 -2608 -4787
rect -2889 -4817 -2859 -4816
rect -2889 -4821 -2858 -4817
rect -3090 -4833 -3086 -4823
rect -2889 -4833 -2884 -4821
rect -2867 -4822 -2858 -4821
rect -2835 -4818 -2831 -4811
rect -2786 -4818 -2782 -4808
rect -2619 -4791 -2608 -4788
rect -2619 -4801 -2616 -4791
rect -2601 -4792 -2597 -4779
rect -2619 -4814 -2616 -4806
rect -2609 -4807 -2605 -4802
rect -2591 -4807 -2590 -4803
rect -2619 -4818 -2609 -4814
rect -2835 -4823 -2794 -4818
rect -2786 -4823 -2723 -4818
rect -2835 -4826 -2831 -4823
rect -2786 -4826 -2782 -4823
rect -3141 -4837 -3129 -4833
rect -3168 -4854 -3162 -4837
rect -3168 -4859 -3155 -4854
rect -3149 -4859 -3143 -4854
rect -3133 -4862 -3129 -4837
rect -3116 -4838 -3098 -4833
rect -3090 -4838 -2910 -4833
rect -2904 -4838 -2884 -4833
rect -2850 -4830 -2813 -4826
rect -2850 -4836 -2846 -4830
rect -2817 -4836 -2813 -4830
rect -3090 -4850 -3086 -4838
rect -2794 -4846 -2790 -4836
rect -3098 -4867 -3094 -4861
rect -2858 -4853 -2854 -4846
rect -2825 -4853 -2821 -4846
rect -2802 -4847 -2775 -4846
rect -2802 -4851 -2801 -4847
rect -2797 -4851 -2780 -4847
rect -2776 -4851 -2775 -4847
rect -2802 -4852 -2775 -4851
rect -2866 -4854 -2839 -4853
rect -2866 -4858 -2865 -4854
rect -2861 -4858 -2844 -4854
rect -2840 -4858 -2839 -4854
rect -2866 -4859 -2839 -4858
rect -2833 -4854 -2806 -4853
rect -2833 -4858 -2832 -4854
rect -2828 -4858 -2811 -4854
rect -2807 -4858 -2806 -4854
rect -2833 -4859 -2806 -4858
rect -2728 -4865 -2723 -4823
rect -2626 -4835 -2622 -4829
rect -2601 -4835 -2597 -4834
rect -2626 -4838 -2597 -4835
rect -2601 -4841 -2597 -4838
rect -2591 -4841 -2587 -4834
rect -2630 -4845 -2608 -4841
rect -2601 -4845 -2587 -4841
rect -2630 -4846 -2613 -4845
rect -2630 -4865 -2625 -4846
rect -3106 -4868 -3079 -4867
rect -3106 -4872 -3105 -4868
rect -3101 -4872 -3084 -4868
rect -3080 -4872 -3079 -4868
rect -3106 -4873 -3079 -4872
rect -3141 -4888 -3137 -4882
rect -3149 -4889 -3122 -4888
rect -3149 -4893 -3148 -4889
rect -3144 -4893 -3127 -4889
rect -3123 -4893 -3122 -4889
rect -3149 -4894 -3122 -4893
rect -2999 -4921 -2994 -4867
rect -2937 -4875 -2933 -4865
rect -2728 -4870 -2625 -4865
rect -2616 -4865 -2613 -4846
rect -2601 -4846 -2597 -4845
rect -2591 -4846 -2587 -4845
rect -2583 -4841 -2579 -4834
rect -2583 -4845 -2567 -4841
rect -2583 -4846 -2579 -4845
rect -2609 -4857 -2605 -4856
rect -2592 -4861 -2584 -4857
rect -2580 -4861 -2578 -4857
rect -2570 -4865 -2567 -4845
rect -2616 -4868 -2567 -4865
rect -2947 -4907 -2936 -4903
rect -2963 -4912 -2944 -4907
rect -2929 -4908 -2925 -4895
rect -2963 -4921 -2958 -4912
rect -2999 -4926 -2958 -4921
rect -2947 -4917 -2944 -4912
rect -2947 -4930 -2944 -4922
rect -2937 -4923 -2933 -4918
rect -2919 -4923 -2918 -4919
rect -2947 -4934 -2937 -4930
rect -2929 -4957 -2925 -4950
rect -2919 -4957 -2915 -4950
rect -2944 -4961 -2936 -4957
rect -2929 -4961 -2915 -4957
rect -2944 -4964 -2941 -4961
rect -2929 -4962 -2925 -4961
rect -2919 -4962 -2915 -4961
rect -2911 -4957 -2907 -4950
rect -2911 -4961 -2895 -4957
rect -2911 -4962 -2907 -4961
rect -2944 -4981 -2941 -4969
rect -2937 -4973 -2933 -4972
rect -2920 -4977 -2912 -4973
rect -2908 -4977 -2906 -4973
rect -2898 -4981 -2895 -4961
rect -2944 -4984 -2895 -4981
<< m2contact >>
rect 1815 368 1821 373
rect 1785 286 1791 291
rect -2970 -2108 -2961 -2103
rect -3184 -2183 -3175 -2178
rect -2897 -2229 -2891 -2224
rect -3115 -2390 -3109 -2385
rect -3158 -2456 -3152 -2451
rect -3145 -2472 -3139 -2467
rect -3073 -2451 -3067 -2446
rect -2927 -2311 -2921 -2306
rect -2752 -2267 -2746 -2262
rect -2559 -2283 -2553 -2278
rect -2782 -2349 -2776 -2344
rect -2710 -2328 -2704 -2323
rect -2413 -2281 -2407 -2276
rect -2269 -2285 -2263 -2280
rect -2325 -2311 -2317 -2306
rect -2602 -2365 -2594 -2359
rect -2589 -2365 -2583 -2360
rect -2443 -2363 -2437 -2358
rect -2114 -2287 -2108 -2282
rect -2331 -2398 -2326 -2393
rect -2299 -2367 -2293 -2362
rect -1979 -2295 -1973 -2290
rect -2144 -2369 -2138 -2364
rect -1870 -2322 -1864 -2317
rect -2022 -2377 -2016 -2372
rect -2009 -2377 -2003 -2372
rect -1877 -2373 -1870 -2368
rect -1574 -2411 -1569 -2406
rect -1558 -2483 -1553 -2478
rect -1391 -2560 -1385 -2555
rect -2662 -2949 -2657 -2944
rect -2373 -2843 -2368 -2838
rect -3122 -3305 -3116 -3300
rect -2889 -3044 -2883 -3039
rect -2949 -3069 -2937 -3064
rect -2662 -2979 -2657 -2974
rect -2720 -3043 -2714 -3038
rect -2768 -3067 -2763 -3061
rect -2556 -3041 -2550 -3036
rect -2416 -3043 -2410 -3038
rect -2476 -3067 -2471 -3062
rect -2932 -3126 -2923 -3120
rect -2919 -3126 -2913 -3121
rect -2750 -3125 -2744 -3120
rect -2586 -3123 -2580 -3118
rect -2265 -3056 -2259 -3051
rect -2456 -3126 -2450 -3120
rect -2446 -3125 -2440 -3120
rect -2350 -3104 -2343 -3099
rect -2295 -3138 -2289 -3133
rect -2020 -3119 -2010 -3114
rect -2102 -3260 -2096 -3255
rect -2543 -3337 -2538 -3332
rect -2168 -3335 -2163 -3330
rect -2132 -3342 -2126 -3337
rect -3152 -3387 -3146 -3382
rect -1752 -3489 -1745 -3484
rect -1487 -3456 -1482 -3451
rect -1500 -3527 -1495 -3522
rect -1487 -3527 -1482 -3522
rect -1468 -3527 -1463 -3522
rect -3128 -4154 -3122 -4149
rect -2868 -3817 -2862 -3812
rect -2939 -3842 -2934 -3837
rect -2930 -3842 -2925 -3837
rect -2962 -3883 -2953 -3876
rect -2898 -3899 -2892 -3894
rect -2867 -4022 -2861 -4017
rect -2923 -4046 -2918 -4041
rect -2910 -4104 -2904 -4099
rect -2897 -4104 -2891 -4099
rect -2633 -4093 -2623 -4088
rect -2427 -4068 -2422 -4063
rect -2405 -4067 -2400 -4062
rect -2992 -4197 -2987 -4192
rect -2418 -4138 -2413 -4133
rect -2405 -4138 -2400 -4133
rect -2386 -4138 -2381 -4133
rect 720 -4167 725 -4162
rect -3158 -4236 -3152 -4231
rect -2992 -4231 -2987 -4226
rect 707 -4238 712 -4233
rect 720 -4238 725 -4233
rect 739 -4238 744 -4233
rect -2963 -4380 -2954 -4373
rect -2886 -4380 -2878 -4373
rect -2956 -4597 -2950 -4592
rect -3008 -4621 -3003 -4616
rect -3125 -4777 -3119 -4772
rect -3031 -4821 -3026 -4816
rect -2986 -4679 -2980 -4674
rect -2885 -4770 -2878 -4765
rect -2999 -4822 -2994 -4812
rect -2597 -4791 -2592 -4786
rect -3155 -4859 -3149 -4854
rect -2910 -4838 -2904 -4833
rect -2999 -4867 -2994 -4852
rect -2610 -4862 -2605 -4857
rect -2597 -4862 -2592 -4857
rect -2578 -4862 -2573 -4857
rect -2925 -4907 -2920 -4902
rect -2946 -4969 -2941 -4964
rect -2938 -4978 -2933 -4973
rect -2925 -4978 -2920 -4973
rect -2906 -4978 -2901 -4973
<< metal2 >>
rect 1815 303 1821 368
rect 1785 296 1821 303
rect 1785 291 1791 296
rect -2993 -2041 -1424 -2036
rect -3198 -2183 -3184 -2178
rect -3198 -2184 -3175 -2183
rect -3198 -2451 -3192 -2184
rect -3198 -2456 -3158 -2451
rect -3115 -2455 -3109 -2390
rect -2993 -2446 -2988 -2041
rect -2970 -2113 -2961 -2108
rect -3067 -2451 -2988 -2446
rect -3198 -2457 -3152 -2456
rect -3158 -2459 -3152 -2457
rect -3145 -2462 -3109 -2455
rect -3145 -2467 -3139 -2462
rect -2966 -2838 -2961 -2113
rect -2697 -2146 -1894 -2141
rect -2897 -2294 -2891 -2229
rect -2927 -2301 -2891 -2294
rect -2927 -2306 -2921 -2301
rect -2752 -2332 -2746 -2267
rect -2697 -2323 -2692 -2146
rect -2053 -2176 -1913 -2171
rect -2704 -2328 -2692 -2323
rect -2782 -2339 -2746 -2332
rect -2782 -2344 -2776 -2339
rect -2559 -2348 -2553 -2283
rect -2413 -2346 -2407 -2281
rect -2589 -2355 -2553 -2348
rect -2443 -2353 -2407 -2346
rect -2343 -2311 -2325 -2306
rect -2655 -2365 -2602 -2359
rect -2589 -2360 -2583 -2355
rect -2443 -2358 -2437 -2353
rect -2655 -2366 -2594 -2365
rect -2655 -2753 -2648 -2366
rect -2343 -2438 -2338 -2311
rect -2269 -2350 -2263 -2285
rect -2299 -2357 -2263 -2350
rect -2114 -2352 -2108 -2287
rect -2299 -2362 -2293 -2357
rect -2144 -2359 -2108 -2352
rect -2144 -2364 -2138 -2359
rect -2331 -2424 -2326 -2398
rect -2053 -2424 -2048 -2176
rect -1979 -2360 -1973 -2295
rect -2009 -2367 -1973 -2360
rect -2331 -2429 -2048 -2424
rect -2036 -2372 -2016 -2371
rect -2036 -2377 -2022 -2372
rect -2009 -2372 -2003 -2367
rect -1918 -2368 -1913 -2176
rect -1899 -2317 -1894 -2146
rect -1899 -2322 -1870 -2317
rect -1918 -2373 -1877 -2368
rect -2036 -2378 -2016 -2377
rect -2343 -2443 -2192 -2438
rect -2655 -2760 -2343 -2753
rect -2966 -2843 -2373 -2838
rect -2787 -2940 -2471 -2935
rect -2949 -3103 -2945 -3069
rect -2952 -3105 -2945 -3103
rect -2952 -3107 -2946 -3105
rect -3021 -3113 -2946 -3107
rect -2889 -3109 -2883 -3044
rect -2787 -3074 -2782 -2940
rect -2662 -2974 -2657 -2949
rect -2768 -3074 -2763 -3067
rect -2787 -3079 -2763 -3074
rect -3122 -3370 -3116 -3305
rect -3152 -3377 -3116 -3370
rect -3152 -3382 -3146 -3377
rect -3128 -4219 -3122 -4154
rect -3158 -4226 -3122 -4219
rect -3158 -4231 -3152 -4226
rect -3125 -4842 -3119 -4777
rect -3155 -4849 -3119 -4842
rect -3155 -4854 -3149 -4849
rect -3031 -4969 -3026 -4821
rect -3021 -4825 -3015 -3113
rect -2919 -3116 -2883 -3109
rect -2949 -3126 -2932 -3120
rect -2919 -3121 -2913 -3116
rect -2949 -3127 -2941 -3126
rect -3011 -3883 -2962 -3876
rect -3011 -4373 -3005 -3883
rect -2992 -4226 -2987 -4197
rect -3011 -4380 -2963 -4373
rect -2949 -4471 -2945 -3127
rect -2768 -3710 -2763 -3079
rect -2720 -3108 -2714 -3043
rect -2556 -3106 -2550 -3041
rect -2476 -3062 -2471 -2940
rect -2750 -3115 -2714 -3108
rect -2586 -3113 -2550 -3106
rect -2416 -3108 -2410 -3043
rect -2350 -3099 -2343 -2760
rect -2750 -3120 -2744 -3115
rect -2586 -3118 -2580 -3113
rect -2446 -3115 -2410 -3108
rect -2446 -3120 -2440 -3115
rect -2265 -3121 -2259 -3056
rect -2456 -3171 -2450 -3126
rect -2295 -3128 -2259 -3121
rect -2295 -3133 -2289 -3128
rect -2197 -3132 -2192 -2443
rect -2036 -2628 -2029 -2378
rect -1574 -2478 -1569 -2411
rect -1574 -2483 -1558 -2478
rect -1429 -2555 -1424 -2041
rect -1429 -2560 -1391 -2555
rect -2036 -2635 -2002 -2628
rect -2009 -2926 -2002 -2635
rect -2009 -2933 -1745 -2926
rect -2203 -3137 -2192 -3132
rect -2168 -3114 -2015 -3111
rect -2168 -3116 -2020 -3114
rect -2930 -3715 -2763 -3710
rect -2756 -3177 -2450 -3171
rect -2930 -3837 -2925 -3715
rect -2756 -3725 -2750 -3177
rect -2203 -3277 -2198 -3137
rect -2805 -3731 -2750 -3725
rect -2629 -3282 -2198 -3277
rect -2939 -4041 -2934 -3842
rect -2868 -3882 -2862 -3817
rect -2898 -3889 -2862 -3882
rect -2898 -3894 -2892 -3889
rect -2939 -4046 -2923 -4041
rect -2867 -4087 -2861 -4022
rect -2897 -4094 -2861 -4087
rect -2897 -4099 -2891 -4094
rect -3008 -4475 -2945 -4471
rect -2910 -4156 -2904 -4104
rect -2805 -4156 -2799 -3731
rect -2629 -4088 -2624 -3282
rect -2168 -3330 -2163 -3116
rect -2027 -3119 -2020 -3116
rect -2102 -3325 -2096 -3260
rect -2168 -3336 -2163 -3335
rect -2132 -3332 -2096 -3325
rect -2543 -3910 -2538 -3337
rect -2132 -3337 -2126 -3332
rect -1752 -3484 -1745 -2933
rect -1482 -3455 -1464 -3452
rect -1467 -3522 -1464 -3455
rect -1495 -3526 -1487 -3522
rect -2543 -3915 -2484 -3910
rect -2489 -4040 -2484 -3915
rect -2489 -4045 -2446 -4040
rect -2451 -4063 -2446 -4045
rect -2451 -4068 -2427 -4063
rect -2400 -4066 -2382 -4063
rect -2385 -4133 -2382 -4066
rect -2413 -4137 -2405 -4133
rect -2910 -4162 -2799 -4156
rect -3008 -4616 -3004 -4475
rect -2956 -4662 -2950 -4597
rect -2986 -4669 -2950 -4662
rect -2986 -4674 -2980 -4669
rect -2999 -4825 -2994 -4822
rect -3021 -4830 -2994 -4825
rect -2999 -4852 -2994 -4830
rect -2910 -4833 -2904 -4162
rect 725 -4166 743 -4163
rect 740 -4233 743 -4166
rect 712 -4237 720 -4233
rect -2885 -4765 -2878 -4380
rect -2592 -4790 -2574 -4787
rect -2910 -4839 -2904 -4838
rect -2577 -4857 -2574 -4790
rect -2605 -4861 -2597 -4857
rect -2920 -4906 -2902 -4903
rect -2977 -4969 -2946 -4964
rect -3031 -4974 -2972 -4969
rect -2905 -4973 -2902 -4906
rect -2933 -4977 -2925 -4973
<< m123contact >>
rect -1509 -3471 -1504 -3466
rect -1486 -3472 -1481 -3467
rect -2427 -4082 -2422 -4077
rect -2404 -4083 -2399 -4078
rect 698 -4182 703 -4177
rect 721 -4183 726 -4178
rect -2619 -4806 -2614 -4801
rect -2596 -4807 -2591 -4802
rect -2947 -4922 -2942 -4917
rect -2924 -4923 -2919 -4918
<< metal3 >>
rect -1504 -3471 -1486 -3467
rect -2422 -4082 -2404 -4078
rect 703 -4182 721 -4178
rect -2614 -4806 -2596 -4802
rect -2942 -4922 -2924 -4918
<< labels >>
rlabel metal1 2111 321 2111 321 3 gnd
rlabel metal1 2197 321 2197 321 7 vdd
rlabel metal1 2197 270 2197 270 7 vdd
rlabel metal1 2111 270 2111 270 3 gnd
rlabel metal1 2261 342 2261 342 5 vdd
rlabel metal1 2261 269 2261 269 1 gnd
rlabel metal1 2464 159 2464 159 1 gnd
rlabel metal1 2464 232 2464 232 5 vdd
rlabel metal1 2415 280 2415 280 5 vdd
rlabel metal1 2400 152 2400 152 1 gnd
rlabel metal1 2433 152 2433 152 1 gnd
rlabel metal1 1847 275 1847 275 1 gnd
rlabel metal1 1847 371 1847 371 5 vdd
rlabel metal1 1812 441 1812 441 5 vdd
rlabel metal1 1785 441 1785 441 5 vdd
rlabel metal1 1804 254 1804 254 1 gnd
rlabel metal1 -3197 -4533 -3197 -4533 3 gnd
rlabel metal1 -3111 -4533 -3111 -4533 7 vdd
rlabel metal1 -3111 -4584 -3111 -4584 7 vdd
rlabel metal1 -3197 -4584 -3197 -4584 3 gnd
rlabel metal1 -3047 -4512 -3047 -4512 5 vdd
rlabel metal1 -3047 -4585 -3047 -4585 1 gnd
rlabel metal1 -3175 -3771 -3175 -3771 3 gnd
rlabel metal1 -3089 -3771 -3089 -3771 7 vdd
rlabel metal1 -3089 -3822 -3089 -3822 7 vdd
rlabel metal1 -3175 -3822 -3175 -3822 3 gnd
rlabel metal1 -3025 -3750 -3025 -3750 5 vdd
rlabel metal1 -3025 -3823 -3025 -3823 1 gnd
rlabel metal1 -3175 -3003 -3175 -3003 3 gnd
rlabel metal1 -3089 -3003 -3089 -3003 7 vdd
rlabel metal1 -3089 -3054 -3089 -3054 7 vdd
rlabel metal1 -3175 -3054 -3175 -3054 3 gnd
rlabel metal1 -3025 -2982 -3025 -2982 5 vdd
rlabel metal1 -3025 -3055 -3025 -3055 1 gnd
rlabel metal1 -3181 -2152 -3181 -2152 3 gnd
rlabel metal1 -3095 -2152 -3095 -2152 7 vdd
rlabel metal1 -3095 -2203 -3095 -2203 7 vdd
rlabel metal1 -3181 -2203 -3181 -2203 3 gnd
rlabel metal1 -3031 -2131 -3031 -2131 5 vdd
rlabel metal1 -3031 -2204 -3031 -2204 1 gnd
rlabel metal1 -3133 -3419 -3133 -3419 1 gnd
rlabel metal1 -3152 -3232 -3152 -3232 5 vdd
rlabel metal1 -3125 -3232 -3125 -3232 5 vdd
rlabel metal1 -3090 -3302 -3090 -3302 5 vdd
rlabel metal1 -3090 -3398 -3090 -3398 1 gnd
rlabel metal1 -3139 -4268 -3139 -4268 1 gnd
rlabel metal1 -3158 -4081 -3158 -4081 5 vdd
rlabel metal1 -3131 -4081 -3131 -4081 5 vdd
rlabel metal1 -3096 -4151 -3096 -4151 5 vdd
rlabel metal1 -3096 -4247 -3096 -4247 1 gnd
rlabel metal1 -3017 -2175 -3017 -2175 1 p3
rlabel metal1 -3083 -2483 -3083 -2483 1 gnd
rlabel metal1 -3083 -2387 -3083 -2387 5 vdd
rlabel metal1 -3118 -2317 -3118 -2317 5 vdd
rlabel metal1 -3145 -2317 -3145 -2317 5 vdd
rlabel metal1 -3126 -2504 -3126 -2504 1 gnd
rlabel metal1 -3136 -4891 -3136 -4891 1 gnd
rlabel metal1 -3155 -4704 -3155 -4704 5 vdd
rlabel metal1 -3128 -4704 -3128 -4704 5 vdd
rlabel metal1 -3093 -4774 -3093 -4774 5 vdd
rlabel metal1 -3093 -4870 -3093 -4870 1 gnd
rlabel metal1 -3033 -4556 -3033 -4556 1 p0
rlabel metal1 -3081 -4835 -3081 -4835 1 g0
rlabel metal1 -2967 -4711 -2967 -4711 1 gnd
rlabel metal1 -2986 -4524 -2986 -4524 5 vdd
rlabel metal1 -2959 -4524 -2959 -4524 5 vdd
rlabel metal1 -2924 -4594 -2924 -4594 5 vdd
rlabel metal1 -2924 -4690 -2924 -4690 1 gnd
rlabel metal1 -2996 -4913 -2996 -4913 1 c0
rlabel metal1 -2820 -4856 -2820 -4856 1 gnd
rlabel metal1 -2853 -4856 -2853 -4856 1 gnd
rlabel metal1 -2838 -4728 -2838 -4728 5 vdd
rlabel metal1 -2789 -4776 -2789 -4776 5 vdd
rlabel metal1 -2789 -4849 -2789 -4849 1 gnd
rlabel metal1 -2776 -4820 -2776 -4820 1 c1
rlabel metal1 -2879 -3931 -2879 -3931 1 gnd
rlabel metal1 -2898 -3744 -2898 -3744 5 vdd
rlabel metal1 -2871 -3744 -2871 -3744 5 vdd
rlabel metal1 -2836 -3814 -2836 -3814 5 vdd
rlabel metal1 -2836 -3910 -2836 -3910 1 gnd
rlabel metal1 -2878 -4136 -2878 -4136 1 gnd
rlabel metal1 -2897 -3949 -2897 -3949 5 vdd
rlabel metal1 -2870 -3949 -2870 -3949 5 vdd
rlabel metal1 -2835 -4019 -2835 -4019 5 vdd
rlabel metal1 -2835 -4115 -2835 -4115 1 gnd
rlabel metal1 -3084 -4212 -3084 -4212 1 g1
rlabel metal1 -2823 -3875 -2823 -3875 1 0c2
rlabel metal1 -2821 -4081 -2821 -4081 1 1c2
rlabel metal1 -2683 -4006 -2683 -4006 1 gnd
rlabel metal1 -2683 -3933 -2683 -3933 5 vdd
rlabel metal1 -2732 -3885 -2732 -3885 5 vdd
rlabel metal1 -2747 -4013 -2747 -4013 1 gnd
rlabel metal1 -2714 -4013 -2714 -4013 1 gnd
rlabel metal1 -2537 -4119 -2537 -4119 1 gnd
rlabel metal1 -2537 -4046 -2537 -4046 5 vdd
rlabel metal1 -2586 -3998 -2586 -3998 5 vdd
rlabel metal1 -2601 -4126 -2601 -4126 1 gnd
rlabel metal1 -2568 -4126 -2568 -4126 1 gnd
rlabel metal1 -2645 -3978 -2645 -3978 1 2c2
rlabel metal1 -2523 -4090 -2523 -4090 1 c2
rlabel metal1 -2857 -3137 -2857 -3137 1 gnd
rlabel metal1 -2857 -3041 -2857 -3041 5 vdd
rlabel metal1 -2892 -2971 -2892 -2971 5 vdd
rlabel metal1 -2919 -2971 -2919 -2971 5 vdd
rlabel metal1 -2900 -3158 -2900 -3158 1 gnd
rlabel metal1 -2731 -3157 -2731 -3157 1 gnd
rlabel metal1 -2750 -2970 -2750 -2970 5 vdd
rlabel metal1 -2723 -2970 -2723 -2970 5 vdd
rlabel metal1 -2688 -3040 -2688 -3040 5 vdd
rlabel metal1 -2688 -3136 -2688 -3136 1 gnd
rlabel metal1 -2567 -3155 -2567 -3155 1 gnd
rlabel metal1 -2586 -2968 -2586 -2968 5 vdd
rlabel metal1 -2559 -2968 -2559 -2968 5 vdd
rlabel metal1 -2524 -3038 -2524 -3038 5 vdd
rlabel metal1 -2524 -3134 -2524 -3134 1 gnd
rlabel metal1 -3012 -3027 -3012 -3027 1 p2
rlabel metal1 -3076 -3364 -3076 -3364 1 g2
rlabel metal1 -2827 -3102 -2827 -3102 1 0c3
rlabel metal1 -2674 -3102 -2674 -3102 1 1c3
rlabel metal1 -2510 -3099 -2510 -3099 1 2c3
rlabel metal1 -2384 -3136 -2384 -3136 1 gnd
rlabel metal1 -2384 -3040 -2384 -3040 5 vdd
rlabel metal1 -2419 -2970 -2419 -2970 5 vdd
rlabel metal1 -2446 -2970 -2446 -2970 5 vdd
rlabel metal1 -2427 -3157 -2427 -3157 1 gnd
rlabel metal1 -2070 -3353 -2070 -3353 1 gnd
rlabel metal1 -2070 -3257 -2070 -3257 5 vdd
rlabel metal1 -2105 -3187 -2105 -3187 5 vdd
rlabel metal1 -2132 -3187 -2132 -3187 5 vdd
rlabel metal1 -2113 -3374 -2113 -3374 1 gnd
rlabel metal1 -2369 -3102 -2369 -3102 1 3c3
rlabel metal1 -2056 -3319 -2056 -3319 1 5c3
rlabel metal1 -1967 -3153 -1967 -3153 1 gnd
rlabel metal1 -2000 -3153 -2000 -3153 1 gnd
rlabel metal1 -1985 -3025 -1985 -3025 5 vdd
rlabel metal1 -1936 -3073 -1936 -3073 5 vdd
rlabel metal1 -1936 -3146 -1936 -3146 1 gnd
rlabel metal1 -1802 -3356 -1802 -3356 1 gnd
rlabel metal1 -1802 -3283 -1802 -3283 5 vdd
rlabel metal1 -1851 -3235 -1851 -3235 5 vdd
rlabel metal1 -1866 -3363 -1866 -3363 1 gnd
rlabel metal1 -1833 -3363 -1833 -3363 1 gnd
rlabel metal1 -1655 -3516 -1655 -3516 1 gnd
rlabel metal1 -1655 -3443 -1655 -3443 5 vdd
rlabel metal1 -1704 -3395 -1704 -3395 5 vdd
rlabel metal1 -1719 -3523 -1719 -3523 1 gnd
rlabel metal1 -1686 -3523 -1686 -3523 1 gnd
rlabel metal1 -1924 -3117 -1924 -3117 1 6c3
rlabel metal1 -1787 -3328 -1787 -3328 1 7c3
rlabel metal1 -1641 -3487 -1641 -3487 1 c3
rlabel metal1 -2865 -2322 -2865 -2322 1 gnd
rlabel metal1 -2865 -2226 -2865 -2226 5 vdd
rlabel metal1 -2900 -2156 -2900 -2156 5 vdd
rlabel metal1 -2927 -2156 -2927 -2156 5 vdd
rlabel metal1 -2908 -2343 -2908 -2343 1 gnd
rlabel metal1 -2852 -2287 -2852 -2287 1 2c4
rlabel metal1 -2763 -2381 -2763 -2381 1 gnd
rlabel metal1 -2782 -2194 -2782 -2194 5 vdd
rlabel metal1 -2755 -2194 -2755 -2194 5 vdd
rlabel metal1 -2720 -2264 -2720 -2264 5 vdd
rlabel metal1 -2720 -2360 -2720 -2360 1 gnd
rlabel m2contact -2706 -2326 -2706 -2326 1 3c3
rlabel metal1 -2527 -2376 -2527 -2376 1 gnd
rlabel metal1 -2527 -2280 -2527 -2280 5 vdd
rlabel metal1 -2562 -2210 -2562 -2210 5 vdd
rlabel metal1 -2589 -2210 -2589 -2210 5 vdd
rlabel metal1 -2570 -2397 -2570 -2397 1 gnd
rlabel metal1 -2381 -2374 -2381 -2374 1 gnd
rlabel metal1 -2381 -2278 -2381 -2278 5 vdd
rlabel metal1 -2416 -2208 -2416 -2208 5 vdd
rlabel metal1 -2443 -2208 -2443 -2208 5 vdd
rlabel metal1 -2424 -2395 -2424 -2395 1 gnd
rlabel metal1 -2514 -2341 -2514 -2341 1 5c4
rlabel metal1 -2367 -2339 -2367 -2339 1 6c4
rlabel metal1 -2237 -2378 -2237 -2378 1 gnd
rlabel metal1 -2237 -2282 -2237 -2282 5 vdd
rlabel metal1 -2272 -2212 -2272 -2212 5 vdd
rlabel metal1 -2299 -2212 -2299 -2212 5 vdd
rlabel metal1 -2280 -2399 -2280 -2399 1 gnd
rlabel metal1 -2082 -2380 -2082 -2380 1 gnd
rlabel metal1 -2082 -2284 -2082 -2284 5 vdd
rlabel metal1 -2117 -2214 -2117 -2214 5 vdd
rlabel metal1 -2144 -2214 -2144 -2214 5 vdd
rlabel metal1 -2125 -2401 -2125 -2401 1 gnd
rlabel metal1 -2233 -3149 -2233 -3149 1 gnd
rlabel metal1 -2233 -3053 -2233 -3053 5 vdd
rlabel metal1 -2268 -2983 -2268 -2983 5 vdd
rlabel metal1 -2295 -2983 -2295 -2983 5 vdd
rlabel metal1 -2276 -3170 -2276 -3170 1 gnd
rlabel metal1 -2220 -3115 -2220 -3115 1 4c3
rlabel metal1 -2223 -2343 -2223 -2343 1 7c4
rlabel metal1 -2068 -2346 -2068 -2346 1 8c4
rlabel metal1 -1947 -2388 -1947 -2388 1 gnd
rlabel metal1 -1947 -2292 -1947 -2292 5 vdd
rlabel metal1 -1982 -2222 -1982 -2222 5 vdd
rlabel metal1 -2009 -2222 -2009 -2222 5 vdd
rlabel metal1 -1990 -2409 -1990 -2409 1 gnd
rlabel metal1 -1933 -2353 -1933 -2353 1 9c4
rlabel metal1 -1799 -2399 -1799 -2399 1 gnd
rlabel metal1 -1799 -2326 -1799 -2326 5 vdd
rlabel metal1 -1848 -2278 -1848 -2278 5 vdd
rlabel metal1 -1863 -2406 -1863 -2406 1 gnd
rlabel metal1 -1830 -2406 -1830 -2406 1 gnd
rlabel metal1 -1668 -2462 -1668 -2462 1 gnd
rlabel metal1 -1701 -2462 -1701 -2462 1 gnd
rlabel metal1 -1686 -2334 -1686 -2334 5 vdd
rlabel metal1 -1637 -2382 -1637 -2382 5 vdd
rlabel metal1 -1637 -2455 -1637 -2455 1 gnd
rlabel metal1 -1510 -2518 -1510 -2518 1 gnd
rlabel metal1 -1543 -2518 -1543 -2518 1 gnd
rlabel metal1 -1528 -2390 -1528 -2390 5 vdd
rlabel metal1 -1479 -2438 -1479 -2438 5 vdd
rlabel metal1 -1479 -2511 -1479 -2511 1 gnd
rlabel metal1 -1344 -2594 -1344 -2594 1 gnd
rlabel metal1 -1377 -2594 -1377 -2594 1 gnd
rlabel metal1 -1362 -2466 -1362 -2466 5 vdd
rlabel metal1 -1313 -2514 -1313 -2514 5 vdd
rlabel metal1 -1313 -2587 -1313 -2587 1 gnd
rlabel metal1 -1785 -2371 -1785 -2371 1 10c4
rlabel metal1 -1624 -2426 -1624 -2426 1 11c4
rlabel metal1 -1466 -2483 -1466 -2483 1 12c4
rlabel m2contact -3069 -2448 -3069 -2448 1 g3
rlabel metal1 -1300 -2559 -1300 -2559 1 c4
rlabel metal1 -3179 -4799 -3179 -4799 1 a0
rlabel metal1 -3166 -4839 -3166 -4839 1 b0
rlabel metal1 -3196 -4515 -3196 -4515 1 a0
rlabel metal1 -3196 -4562 -3196 -4562 1 b0
rlabel metal1 -3168 -4218 -3168 -4218 1 b1
rlabel metal1 -3174 -4174 -3174 -4174 1 a1
rlabel metal1 -3176 -3800 -3176 -3800 1 b1
rlabel metal1 -3174 -3753 -3174 -3753 1 a1
rlabel metal1 -3162 -3369 -3162 -3369 1 b2
rlabel metal1 -3167 -3320 -3167 -3320 1 a2
rlabel metal1 -3175 -3031 -3175 -3031 1 b2
rlabel metal1 -3172 -2984 -3172 -2984 1 a2
rlabel metal1 -3175 -2134 -3175 -2134 1 a3
rlabel metal2 -3196 -2182 -3196 -2182 1 b3
rlabel metal1 703 -4166 705 -4164 3 a
rlabel metal1 703 -4220 705 -4218 1 b
rlabel metal1 709 -4183 711 -4182 1 gnd
rlabel metal1 709 -4128 711 -4126 5 vdd
rlabel metal1 721 -4220 725 -4218 1 out
rlabel metal1 717 -4166 719 -4163 1 a_bar
rlabel metal1 -2608 -4807 -2606 -4806 1 gnd
rlabel metal1 -2600 -4790 -2598 -4787 1 a_bar
rlabel metal1 -2716 -4766 -2716 -4766 1 p1
rlabel metal1 -2624 -4831 -2624 -4831 1 s1
rlabel metal1 -2936 -4923 -2934 -4922 1 gnd
rlabel metal1 -2936 -4868 -2934 -4866 5 vdd
rlabel metal1 -2928 -4906 -2926 -4903 1 a_bar
rlabel metal1 -2416 -4083 -2414 -4082 1 gnd
rlabel metal1 -2416 -4028 -2414 -4026 5 vdd
rlabel metal1 -2408 -4066 -2406 -4063 1 a_bar
rlabel metal1 -1498 -3472 -1496 -3471 1 gnd
rlabel metal1 -1498 -3417 -1496 -3415 5 vdd
rlabel metal1 -1490 -3455 -1488 -3452 1 a_bar
rlabel metal1 -1484 -3509 -1484 -3509 1 s3
rlabel metal1 -2402 -4118 -2402 -4118 1 s2
rlabel metal1 -2922 -4959 -2922 -4959 1 s0
<< end >>
