magic
tech scmos
timestamp 1732103761
<< nwell >>
rect -2926 -538 -2872 -476
rect -2864 -608 -2837 -546
rect -2548 -615 -2496 -588
rect -2450 -620 -2423 -575
rect -2548 -666 -2496 -639
rect -2296 -733 -2269 -637
rect -2247 -730 -2220 -685
rect -2000 -779 -1968 -653
rect -1948 -779 -1916 -653
rect -1896 -717 -1864 -653
rect -1844 -717 -1812 -653
rect -1799 -709 -1735 -645
rect -8323 -3102 -8291 -2976
rect -8271 -3102 -8239 -2976
rect -8219 -3040 -8187 -2976
rect -8167 -3040 -8135 -2976
rect -8122 -3032 -8058 -2968
rect -7840 -3088 -7788 -3061
rect -7742 -3093 -7715 -3048
rect -7840 -3139 -7788 -3112
rect -7638 -3135 -7584 -3073
rect -7576 -3205 -7549 -3143
rect -7493 -3173 -7439 -3111
rect -8309 -3406 -8277 -3280
rect -8257 -3406 -8225 -3280
rect -8205 -3344 -8173 -3280
rect -8153 -3344 -8121 -3280
rect -8108 -3336 -8044 -3272
rect -7856 -3296 -7802 -3234
rect -7431 -3243 -7404 -3181
rect -7300 -3189 -7246 -3127
rect -7154 -3187 -7100 -3125
rect -7010 -3191 -6956 -3129
rect -6855 -3193 -6801 -3131
rect -7238 -3259 -7211 -3197
rect -7092 -3257 -7065 -3195
rect -6948 -3261 -6921 -3199
rect -6720 -3201 -6666 -3139
rect -6793 -3263 -6766 -3201
rect -6658 -3271 -6631 -3209
rect -6559 -3291 -6532 -3195
rect -6510 -3288 -6483 -3243
rect -7794 -3366 -7767 -3304
rect -6397 -3347 -6370 -3251
rect -6348 -3344 -6321 -3299
rect -6239 -3403 -6212 -3307
rect -6190 -3400 -6163 -3355
rect -6073 -3479 -6046 -3383
rect -6024 -3476 -5997 -3431
rect -5923 -3556 -5891 -3430
rect -5871 -3556 -5839 -3430
rect -5819 -3494 -5787 -3430
rect -5767 -3494 -5735 -3430
rect -5722 -3486 -5658 -3422
rect -5553 -3526 -5526 -3464
rect -8254 -4014 -8222 -3888
rect -8202 -4014 -8170 -3888
rect -8150 -3952 -8118 -3888
rect -8098 -3952 -8066 -3888
rect -8053 -3944 -7989 -3880
rect -7834 -3939 -7782 -3912
rect -7736 -3944 -7709 -3899
rect -7630 -3950 -7576 -3888
rect -7461 -3949 -7407 -3887
rect -7297 -3947 -7243 -3885
rect -7157 -3949 -7103 -3887
rect -7834 -3990 -7782 -3963
rect -7568 -4020 -7541 -3958
rect -7399 -4019 -7372 -3957
rect -7235 -4017 -7208 -3955
rect -7095 -4019 -7068 -3957
rect -7006 -3962 -6952 -3900
rect -6944 -4032 -6917 -3970
rect -6696 -4038 -6669 -3942
rect -6647 -4035 -6620 -3990
rect -8237 -4255 -8205 -4129
rect -8185 -4255 -8153 -4129
rect -8133 -4193 -8101 -4129
rect -8081 -4193 -8049 -4129
rect -8036 -4185 -7972 -4121
rect -7863 -4211 -7809 -4149
rect -6843 -4166 -6789 -4104
rect -7801 -4281 -7774 -4219
rect -6781 -4236 -6754 -4174
rect -6562 -4248 -6535 -4152
rect -6513 -4245 -6486 -4200
rect -6415 -4408 -6388 -4312
rect -6366 -4405 -6339 -4360
rect -6203 -4372 -6179 -4340
rect -6203 -4427 -6161 -4395
rect -6090 -4481 -6058 -4355
rect -6038 -4481 -6006 -4355
rect -5986 -4419 -5954 -4355
rect -5934 -4419 -5902 -4355
rect -5889 -4411 -5825 -4347
rect -5729 -4438 -5702 -4376
rect -8248 -4818 -8216 -4692
rect -8196 -4818 -8164 -4692
rect -8144 -4756 -8112 -4692
rect -8092 -4756 -8060 -4692
rect -8047 -4748 -7983 -4684
rect -7834 -4707 -7782 -4680
rect -7736 -4712 -7709 -4667
rect -7609 -4723 -7555 -4661
rect -7834 -4758 -7782 -4731
rect -7547 -4793 -7520 -4731
rect -7608 -4928 -7554 -4866
rect -7443 -4898 -7416 -4802
rect -7394 -4895 -7367 -4850
rect -8235 -5130 -8203 -5004
rect -8183 -5130 -8151 -5004
rect -8131 -5068 -8099 -5004
rect -8079 -5068 -8047 -5004
rect -8034 -5060 -7970 -4996
rect -7546 -4998 -7519 -4936
rect -7869 -5060 -7815 -4998
rect -7297 -5011 -7270 -4915
rect -7248 -5008 -7221 -4963
rect -7121 -4983 -7097 -4951
rect -7121 -5038 -7079 -5006
rect -7807 -5130 -7780 -5068
rect -7009 -5090 -6977 -4964
rect -6957 -5090 -6925 -4964
rect -6905 -5028 -6873 -4964
rect -6853 -5028 -6821 -4964
rect -6808 -5020 -6744 -4956
rect -6695 -5058 -6668 -4996
rect -3996 -5083 -3972 -5051
rect -3996 -5138 -3954 -5106
rect -8248 -5524 -8216 -5398
rect -8196 -5524 -8164 -5398
rect -8144 -5462 -8112 -5398
rect -8092 -5462 -8060 -5398
rect -8047 -5454 -7983 -5390
rect -7856 -5469 -7804 -5442
rect -7758 -5474 -7731 -5429
rect -7856 -5520 -7804 -5493
rect -7697 -5503 -7643 -5441
rect -7635 -5573 -7608 -5511
rect -8245 -5773 -8213 -5647
rect -8193 -5773 -8161 -5647
rect -8141 -5711 -8109 -5647
rect -8089 -5711 -8057 -5647
rect -8044 -5703 -7980 -5639
rect -7866 -5683 -7812 -5621
rect -7804 -5753 -7777 -5691
rect -7549 -5741 -7522 -5645
rect -7500 -5738 -7473 -5693
rect -7313 -5707 -7289 -5675
rect -7313 -5762 -7271 -5730
rect -7193 -5744 -7161 -5618
rect -7141 -5744 -7109 -5618
rect -7089 -5682 -7057 -5618
rect -7037 -5682 -7005 -5618
rect -6992 -5674 -6928 -5610
rect -6831 -5733 -6804 -5671
rect -7641 -5823 -7617 -5791
rect -7641 -5878 -7599 -5846
rect -7870 -6084 -7838 -5958
rect -7818 -6084 -7786 -5958
rect -7766 -6022 -7734 -5958
rect -7714 -6022 -7682 -5958
rect -7669 -6014 -7605 -5950
rect -7470 -5984 -7438 -5858
rect -7418 -5984 -7386 -5858
rect -7366 -5922 -7334 -5858
rect -7314 -5922 -7282 -5858
rect -7269 -5914 -7205 -5850
rect -7132 -5955 -7105 -5893
rect -7556 -6200 -7529 -6138
<< ntransistor >>
rect -2894 -604 -2892 -584
rect -2578 -603 -2568 -601
rect -2473 -615 -2471 -605
rect -2851 -638 -2849 -627
rect -2894 -659 -2892 -639
rect -2473 -648 -2471 -638
rect -2437 -640 -2435 -630
rect -2578 -654 -2568 -652
rect -2234 -750 -2232 -740
rect -2298 -760 -2296 -750
rect -2265 -760 -2263 -750
rect -1784 -740 -1782 -720
rect -1752 -740 -1750 -720
rect -1881 -764 -1879 -744
rect -1829 -764 -1827 -744
rect -1985 -811 -1983 -791
rect -1933 -811 -1931 -791
rect -1881 -811 -1879 -791
rect -1829 -811 -1827 -791
rect -8107 -3063 -8105 -3043
rect -8075 -3063 -8073 -3043
rect -8204 -3087 -8202 -3067
rect -8152 -3087 -8150 -3067
rect -7870 -3076 -7860 -3074
rect -7765 -3088 -7763 -3080
rect -8308 -3134 -8306 -3114
rect -8256 -3134 -8254 -3114
rect -8204 -3134 -8202 -3114
rect -8152 -3134 -8150 -3114
rect -7765 -3121 -7763 -3111
rect -7729 -3113 -7727 -3103
rect -7870 -3127 -7860 -3125
rect -7606 -3201 -7604 -3181
rect -7563 -3235 -7561 -3224
rect -7606 -3256 -7604 -3236
rect -7461 -3239 -7459 -3219
rect -7268 -3255 -7266 -3235
rect -7418 -3273 -7416 -3262
rect -7461 -3294 -7459 -3274
rect -7122 -3253 -7120 -3233
rect -6978 -3257 -6976 -3237
rect -7225 -3289 -7223 -3278
rect -7079 -3287 -7077 -3276
rect -6823 -3259 -6821 -3239
rect -7268 -3310 -7266 -3290
rect -7122 -3308 -7120 -3288
rect -6935 -3291 -6933 -3280
rect -6688 -3267 -6686 -3247
rect -6978 -3312 -6976 -3292
rect -6780 -3293 -6778 -3282
rect -6823 -3314 -6821 -3294
rect -6645 -3301 -6643 -3290
rect -8093 -3367 -8091 -3347
rect -8061 -3367 -8059 -3347
rect -7824 -3362 -7822 -3342
rect -6688 -3322 -6686 -3302
rect -6497 -3308 -6495 -3298
rect -6561 -3318 -6559 -3308
rect -6528 -3318 -6526 -3308
rect -8190 -3391 -8188 -3371
rect -8138 -3391 -8136 -3371
rect -6335 -3364 -6333 -3354
rect -6399 -3374 -6397 -3364
rect -6366 -3374 -6364 -3364
rect -7781 -3396 -7779 -3385
rect -7824 -3417 -7822 -3397
rect -8294 -3438 -8292 -3418
rect -8242 -3438 -8240 -3418
rect -8190 -3438 -8188 -3418
rect -8138 -3438 -8136 -3418
rect -6177 -3420 -6175 -3410
rect -6241 -3430 -6239 -3420
rect -6208 -3430 -6206 -3420
rect -6011 -3496 -6009 -3486
rect -6075 -3506 -6073 -3496
rect -6042 -3506 -6040 -3496
rect -5707 -3517 -5705 -3497
rect -5675 -3517 -5673 -3497
rect -5804 -3541 -5802 -3521
rect -5752 -3541 -5750 -3521
rect -5540 -3556 -5538 -3545
rect -5908 -3588 -5906 -3568
rect -5856 -3588 -5854 -3568
rect -5804 -3588 -5802 -3568
rect -5752 -3588 -5750 -3568
rect -7864 -3927 -7854 -3925
rect -7759 -3939 -7757 -3931
rect -8038 -3975 -8036 -3955
rect -8006 -3975 -8004 -3955
rect -7759 -3972 -7757 -3962
rect -7723 -3964 -7721 -3954
rect -7864 -3978 -7854 -3976
rect -8135 -3999 -8133 -3979
rect -8083 -3999 -8081 -3979
rect -7598 -4016 -7596 -3996
rect -8239 -4046 -8237 -4026
rect -8187 -4046 -8185 -4026
rect -8135 -4046 -8133 -4026
rect -8083 -4046 -8081 -4026
rect -7429 -4015 -7427 -3995
rect -7265 -4013 -7263 -3993
rect -7125 -4015 -7123 -3995
rect -7555 -4050 -7553 -4039
rect -7386 -4049 -7384 -4038
rect -7222 -4047 -7220 -4036
rect -6974 -4028 -6972 -4008
rect -7598 -4071 -7596 -4051
rect -7429 -4070 -7427 -4050
rect -7265 -4068 -7263 -4048
rect -7082 -4049 -7080 -4038
rect -7125 -4070 -7123 -4050
rect -6931 -4062 -6929 -4051
rect -6634 -4055 -6632 -4045
rect -6974 -4083 -6972 -4063
rect -6698 -4065 -6696 -4055
rect -6665 -4065 -6663 -4055
rect -8021 -4216 -8019 -4196
rect -7989 -4216 -7987 -4196
rect -8118 -4240 -8116 -4220
rect -8066 -4240 -8064 -4220
rect -6811 -4232 -6809 -4212
rect -8222 -4287 -8220 -4267
rect -8170 -4287 -8168 -4267
rect -8118 -4287 -8116 -4267
rect -8066 -4287 -8064 -4267
rect -7831 -4277 -7829 -4257
rect -6768 -4266 -6766 -4255
rect -6500 -4265 -6498 -4255
rect -6811 -4287 -6809 -4267
rect -6564 -4275 -6562 -4265
rect -6531 -4275 -6529 -4265
rect -7788 -4311 -7786 -4300
rect -7831 -4332 -7829 -4312
rect -6192 -4389 -6190 -4379
rect -6353 -4425 -6351 -4415
rect -6417 -4435 -6415 -4425
rect -6384 -4435 -6382 -4425
rect -6192 -4443 -6190 -4433
rect -6174 -4443 -6172 -4433
rect -5874 -4442 -5872 -4422
rect -5842 -4442 -5840 -4422
rect -5971 -4466 -5969 -4446
rect -5919 -4466 -5917 -4446
rect -5716 -4468 -5714 -4457
rect -6075 -4513 -6073 -4493
rect -6023 -4513 -6021 -4493
rect -5971 -4513 -5969 -4493
rect -5919 -4513 -5917 -4493
rect -7864 -4695 -7854 -4693
rect -7759 -4707 -7757 -4699
rect -7759 -4740 -7757 -4730
rect -7723 -4732 -7721 -4722
rect -7864 -4746 -7854 -4744
rect -8032 -4779 -8030 -4759
rect -8000 -4779 -7998 -4759
rect -8129 -4803 -8127 -4783
rect -8077 -4803 -8075 -4783
rect -7577 -4789 -7575 -4769
rect -7534 -4823 -7532 -4812
rect -8233 -4850 -8231 -4830
rect -8181 -4850 -8179 -4830
rect -8129 -4850 -8127 -4830
rect -8077 -4850 -8075 -4830
rect -7577 -4844 -7575 -4824
rect -7381 -4915 -7379 -4905
rect -7445 -4925 -7443 -4915
rect -7412 -4925 -7410 -4915
rect -7576 -4994 -7574 -4974
rect -7533 -5028 -7531 -5017
rect -7110 -5000 -7108 -4990
rect -7235 -5028 -7233 -5018
rect -7576 -5049 -7574 -5029
rect -7299 -5038 -7297 -5028
rect -7266 -5038 -7264 -5028
rect -8019 -5091 -8017 -5071
rect -7987 -5091 -7985 -5071
rect -7110 -5054 -7108 -5044
rect -7092 -5054 -7090 -5044
rect -8116 -5115 -8114 -5095
rect -8064 -5115 -8062 -5095
rect -6793 -5051 -6791 -5031
rect -6761 -5051 -6759 -5031
rect -6890 -5075 -6888 -5055
rect -6838 -5075 -6836 -5055
rect -7837 -5126 -7835 -5106
rect -6682 -5088 -6680 -5077
rect -3985 -5100 -3983 -5090
rect -6994 -5122 -6992 -5102
rect -6942 -5122 -6940 -5102
rect -6890 -5122 -6888 -5102
rect -6838 -5122 -6836 -5102
rect -8220 -5162 -8218 -5142
rect -8168 -5162 -8166 -5142
rect -8116 -5162 -8114 -5142
rect -8064 -5162 -8062 -5142
rect -7794 -5160 -7792 -5149
rect -3985 -5154 -3983 -5144
rect -3967 -5154 -3965 -5144
rect -7837 -5181 -7835 -5161
rect -7886 -5457 -7876 -5455
rect -8032 -5485 -8030 -5465
rect -8000 -5485 -7998 -5465
rect -7781 -5469 -7779 -5461
rect -8129 -5509 -8127 -5489
rect -8077 -5509 -8075 -5489
rect -7781 -5502 -7779 -5492
rect -7745 -5494 -7743 -5484
rect -7886 -5508 -7876 -5506
rect -8233 -5556 -8231 -5536
rect -8181 -5556 -8179 -5536
rect -8129 -5556 -8127 -5536
rect -8077 -5556 -8075 -5536
rect -7665 -5569 -7663 -5549
rect -7622 -5603 -7620 -5592
rect -7665 -5624 -7663 -5604
rect -8029 -5734 -8027 -5714
rect -7997 -5734 -7995 -5714
rect -8126 -5758 -8124 -5738
rect -8074 -5758 -8072 -5738
rect -7834 -5749 -7832 -5729
rect -7302 -5724 -7300 -5714
rect -6977 -5705 -6975 -5685
rect -6945 -5705 -6943 -5685
rect -7074 -5729 -7072 -5709
rect -7022 -5729 -7020 -5709
rect -7487 -5758 -7485 -5748
rect -7551 -5768 -7549 -5758
rect -7518 -5768 -7516 -5758
rect -7791 -5783 -7789 -5772
rect -7302 -5778 -7300 -5768
rect -7284 -5778 -7282 -5768
rect -7178 -5776 -7176 -5756
rect -7126 -5776 -7124 -5756
rect -7074 -5776 -7072 -5756
rect -7022 -5776 -7020 -5756
rect -6818 -5763 -6816 -5752
rect -8230 -5805 -8228 -5785
rect -8178 -5805 -8176 -5785
rect -8126 -5805 -8124 -5785
rect -8074 -5805 -8072 -5785
rect -7834 -5804 -7832 -5784
rect -7630 -5840 -7628 -5830
rect -7630 -5894 -7628 -5884
rect -7612 -5894 -7610 -5884
rect -7254 -5945 -7252 -5925
rect -7222 -5945 -7220 -5925
rect -7351 -5969 -7349 -5949
rect -7299 -5969 -7297 -5949
rect -7119 -5985 -7117 -5974
rect -7455 -6016 -7453 -5996
rect -7403 -6016 -7401 -5996
rect -7351 -6016 -7349 -5996
rect -7299 -6016 -7297 -5996
rect -7654 -6045 -7652 -6025
rect -7622 -6045 -7620 -6025
rect -7751 -6069 -7749 -6049
rect -7699 -6069 -7697 -6049
rect -7855 -6116 -7853 -6096
rect -7803 -6116 -7801 -6096
rect -7751 -6116 -7749 -6096
rect -7699 -6116 -7697 -6096
rect -7543 -6230 -7541 -6219
<< ptransistor >>
rect -2913 -530 -2911 -510
rect -2886 -530 -2884 -510
rect -2851 -600 -2849 -560
rect -2540 -603 -2520 -601
rect -2437 -612 -2435 -592
rect -2540 -654 -2520 -652
rect -2283 -678 -2281 -658
rect -2283 -725 -2281 -706
rect -2234 -722 -2232 -702
rect -1985 -708 -1983 -668
rect -1933 -708 -1931 -668
rect -1881 -708 -1879 -668
rect -1829 -708 -1827 -668
rect -1784 -700 -1782 -660
rect -1752 -700 -1750 -660
rect -1985 -770 -1983 -730
rect -1933 -770 -1931 -730
rect -8308 -3031 -8306 -2991
rect -8256 -3031 -8254 -2991
rect -8204 -3031 -8202 -2991
rect -8152 -3031 -8150 -2991
rect -8107 -3023 -8105 -2983
rect -8075 -3023 -8073 -2983
rect -8308 -3093 -8306 -3053
rect -8256 -3093 -8254 -3053
rect -7832 -3076 -7812 -3074
rect -7729 -3085 -7727 -3065
rect -7832 -3127 -7812 -3125
rect -7625 -3127 -7623 -3107
rect -7598 -3127 -7596 -3107
rect -7563 -3197 -7561 -3157
rect -7480 -3165 -7478 -3145
rect -7453 -3165 -7451 -3145
rect -7287 -3181 -7285 -3161
rect -7260 -3181 -7258 -3161
rect -7141 -3179 -7139 -3159
rect -7114 -3179 -7112 -3159
rect -7418 -3235 -7416 -3195
rect -6997 -3183 -6995 -3163
rect -6970 -3183 -6968 -3163
rect -7225 -3251 -7223 -3211
rect -6842 -3185 -6840 -3165
rect -6815 -3185 -6813 -3165
rect -8294 -3335 -8292 -3295
rect -8242 -3335 -8240 -3295
rect -8190 -3335 -8188 -3295
rect -8138 -3335 -8136 -3295
rect -8093 -3327 -8091 -3287
rect -8061 -3327 -8059 -3287
rect -7843 -3288 -7841 -3268
rect -7816 -3288 -7814 -3268
rect -7079 -3249 -7077 -3209
rect -6707 -3193 -6705 -3173
rect -6680 -3193 -6678 -3173
rect -6935 -3253 -6933 -3213
rect -6780 -3255 -6778 -3215
rect -6645 -3263 -6643 -3223
rect -6546 -3236 -6544 -3216
rect -6546 -3283 -6544 -3264
rect -8294 -3397 -8292 -3357
rect -8242 -3397 -8240 -3357
rect -7781 -3358 -7779 -3318
rect -6497 -3280 -6495 -3260
rect -6384 -3292 -6382 -3272
rect -6384 -3339 -6382 -3320
rect -6335 -3336 -6333 -3316
rect -6226 -3348 -6224 -3328
rect -6226 -3395 -6224 -3376
rect -6177 -3392 -6175 -3372
rect -6060 -3424 -6058 -3404
rect -6060 -3471 -6058 -3452
rect -6011 -3468 -6009 -3448
rect -5908 -3485 -5906 -3445
rect -5856 -3485 -5854 -3445
rect -5804 -3485 -5802 -3445
rect -5752 -3485 -5750 -3445
rect -5707 -3477 -5705 -3437
rect -5675 -3477 -5673 -3437
rect -5908 -3547 -5906 -3507
rect -5856 -3547 -5854 -3507
rect -5540 -3518 -5538 -3478
rect -8239 -3943 -8237 -3903
rect -8187 -3943 -8185 -3903
rect -8135 -3943 -8133 -3903
rect -8083 -3943 -8081 -3903
rect -8038 -3935 -8036 -3895
rect -8006 -3935 -8004 -3895
rect -7826 -3927 -7806 -3925
rect -7723 -3936 -7721 -3916
rect -8239 -4005 -8237 -3965
rect -8187 -4005 -8185 -3965
rect -7617 -3942 -7615 -3922
rect -7590 -3942 -7588 -3922
rect -7448 -3941 -7446 -3921
rect -7421 -3941 -7419 -3921
rect -7284 -3939 -7282 -3919
rect -7257 -3939 -7255 -3919
rect -7144 -3941 -7142 -3921
rect -7117 -3941 -7115 -3921
rect -6993 -3954 -6991 -3934
rect -6966 -3954 -6964 -3934
rect -7826 -3978 -7806 -3976
rect -7555 -4012 -7553 -3972
rect -7386 -4011 -7384 -3971
rect -7222 -4009 -7220 -3969
rect -7082 -4011 -7080 -3971
rect -6683 -3983 -6681 -3963
rect -6931 -4024 -6929 -3984
rect -6683 -4030 -6681 -4011
rect -6634 -4027 -6632 -4007
rect -8222 -4184 -8220 -4144
rect -8170 -4184 -8168 -4144
rect -8118 -4184 -8116 -4144
rect -8066 -4184 -8064 -4144
rect -8021 -4176 -8019 -4136
rect -7989 -4176 -7987 -4136
rect -6830 -4158 -6828 -4138
rect -6803 -4158 -6801 -4138
rect -8222 -4246 -8220 -4206
rect -8170 -4246 -8168 -4206
rect -7850 -4203 -7848 -4183
rect -7823 -4203 -7821 -4183
rect -6768 -4228 -6766 -4188
rect -6549 -4193 -6547 -4173
rect -7788 -4273 -7786 -4233
rect -6549 -4240 -6547 -4221
rect -6500 -4237 -6498 -4217
rect -6402 -4353 -6400 -4333
rect -6402 -4400 -6400 -4381
rect -6192 -4366 -6190 -4346
rect -6353 -4397 -6351 -4377
rect -6192 -4421 -6190 -4401
rect -6174 -4421 -6172 -4401
rect -6075 -4410 -6073 -4370
rect -6023 -4410 -6021 -4370
rect -5971 -4410 -5969 -4370
rect -5919 -4410 -5917 -4370
rect -5874 -4402 -5872 -4362
rect -5842 -4402 -5840 -4362
rect -6075 -4472 -6073 -4432
rect -6023 -4472 -6021 -4432
rect -5716 -4430 -5714 -4390
rect -7826 -4695 -7806 -4693
rect -8233 -4747 -8231 -4707
rect -8181 -4747 -8179 -4707
rect -8129 -4747 -8127 -4707
rect -8077 -4747 -8075 -4707
rect -8032 -4739 -8030 -4699
rect -8000 -4739 -7998 -4699
rect -7723 -4704 -7721 -4684
rect -7596 -4715 -7594 -4695
rect -7569 -4715 -7567 -4695
rect -7826 -4746 -7806 -4744
rect -8233 -4809 -8231 -4769
rect -8181 -4809 -8179 -4769
rect -7534 -4785 -7532 -4745
rect -7430 -4843 -7428 -4823
rect -7430 -4890 -7428 -4871
rect -7595 -4920 -7593 -4900
rect -7568 -4920 -7566 -4900
rect -7381 -4887 -7379 -4867
rect -7533 -4990 -7531 -4950
rect -7284 -4956 -7282 -4936
rect -8220 -5059 -8218 -5019
rect -8168 -5059 -8166 -5019
rect -8116 -5059 -8114 -5019
rect -8064 -5059 -8062 -5019
rect -8019 -5051 -8017 -5011
rect -7987 -5051 -7985 -5011
rect -7284 -5003 -7282 -4984
rect -7110 -4977 -7108 -4957
rect -7235 -5000 -7233 -4980
rect -7856 -5052 -7854 -5032
rect -7829 -5052 -7827 -5032
rect -7110 -5032 -7108 -5012
rect -7092 -5032 -7090 -5012
rect -6994 -5019 -6992 -4979
rect -6942 -5019 -6940 -4979
rect -6890 -5019 -6888 -4979
rect -6838 -5019 -6836 -4979
rect -6793 -5011 -6791 -4971
rect -6761 -5011 -6759 -4971
rect -8220 -5121 -8218 -5081
rect -8168 -5121 -8166 -5081
rect -6994 -5081 -6992 -5041
rect -6942 -5081 -6940 -5041
rect -6682 -5050 -6680 -5010
rect -3985 -5077 -3983 -5057
rect -7794 -5122 -7792 -5082
rect -3985 -5132 -3983 -5112
rect -3967 -5132 -3965 -5112
rect -8233 -5453 -8231 -5413
rect -8181 -5453 -8179 -5413
rect -8129 -5453 -8127 -5413
rect -8077 -5453 -8075 -5413
rect -8032 -5445 -8030 -5405
rect -8000 -5445 -7998 -5405
rect -7848 -5457 -7828 -5455
rect -8233 -5515 -8231 -5475
rect -8181 -5515 -8179 -5475
rect -7745 -5466 -7743 -5446
rect -7684 -5495 -7682 -5475
rect -7657 -5495 -7655 -5475
rect -7848 -5508 -7828 -5506
rect -7622 -5565 -7620 -5525
rect -8230 -5702 -8228 -5662
rect -8178 -5702 -8176 -5662
rect -8126 -5702 -8124 -5662
rect -8074 -5702 -8072 -5662
rect -8029 -5694 -8027 -5654
rect -7997 -5694 -7995 -5654
rect -7853 -5675 -7851 -5655
rect -7826 -5675 -7824 -5655
rect -7536 -5686 -7534 -5666
rect -7178 -5673 -7176 -5633
rect -7126 -5673 -7124 -5633
rect -7074 -5673 -7072 -5633
rect -7022 -5673 -7020 -5633
rect -6977 -5665 -6975 -5625
rect -6945 -5665 -6943 -5625
rect -8230 -5764 -8228 -5724
rect -8178 -5764 -8176 -5724
rect -7791 -5745 -7789 -5705
rect -7536 -5733 -7534 -5714
rect -7302 -5701 -7300 -5681
rect -7487 -5730 -7485 -5710
rect -7178 -5735 -7176 -5695
rect -7126 -5735 -7124 -5695
rect -6818 -5725 -6816 -5685
rect -7302 -5756 -7300 -5736
rect -7284 -5756 -7282 -5736
rect -7630 -5817 -7628 -5797
rect -7630 -5872 -7628 -5852
rect -7612 -5872 -7610 -5852
rect -7455 -5913 -7453 -5873
rect -7403 -5913 -7401 -5873
rect -7351 -5913 -7349 -5873
rect -7299 -5913 -7297 -5873
rect -7254 -5905 -7252 -5865
rect -7222 -5905 -7220 -5865
rect -7855 -6013 -7853 -5973
rect -7803 -6013 -7801 -5973
rect -7751 -6013 -7749 -5973
rect -7699 -6013 -7697 -5973
rect -7654 -6005 -7652 -5965
rect -7622 -6005 -7620 -5965
rect -7455 -5975 -7453 -5935
rect -7403 -5975 -7401 -5935
rect -7119 -5947 -7117 -5907
rect -7855 -6075 -7853 -6035
rect -7803 -6075 -7801 -6035
rect -7543 -6192 -7541 -6152
<< ndiffusion >>
rect -2895 -604 -2894 -584
rect -2892 -604 -2891 -584
rect -2578 -601 -2568 -600
rect -2578 -604 -2568 -603
rect -2474 -615 -2473 -605
rect -2471 -615 -2470 -605
rect -2852 -638 -2851 -627
rect -2849 -638 -2848 -627
rect -2895 -659 -2894 -639
rect -2892 -659 -2891 -639
rect -2578 -652 -2568 -651
rect -2474 -648 -2473 -638
rect -2471 -648 -2470 -638
rect -2438 -640 -2437 -630
rect -2435 -640 -2434 -630
rect -2578 -655 -2568 -654
rect -2235 -750 -2234 -740
rect -2232 -750 -2231 -740
rect -2299 -760 -2298 -750
rect -2296 -760 -2295 -750
rect -2266 -760 -2265 -750
rect -2263 -760 -2262 -750
rect -1785 -740 -1784 -720
rect -1782 -740 -1781 -720
rect -1753 -740 -1752 -720
rect -1750 -740 -1749 -720
rect -1882 -764 -1881 -744
rect -1879 -764 -1878 -744
rect -1830 -764 -1829 -744
rect -1827 -764 -1826 -744
rect -1986 -811 -1985 -791
rect -1983 -811 -1982 -791
rect -1934 -811 -1933 -791
rect -1931 -811 -1930 -791
rect -1882 -811 -1881 -791
rect -1879 -811 -1878 -791
rect -1830 -811 -1829 -791
rect -1827 -811 -1826 -791
rect -8108 -3063 -8107 -3043
rect -8105 -3063 -8104 -3043
rect -8076 -3063 -8075 -3043
rect -8073 -3063 -8072 -3043
rect -8205 -3087 -8204 -3067
rect -8202 -3087 -8201 -3067
rect -8153 -3087 -8152 -3067
rect -8150 -3087 -8149 -3067
rect -7870 -3074 -7860 -3073
rect -7870 -3077 -7860 -3076
rect -7766 -3088 -7765 -3080
rect -7763 -3088 -7762 -3080
rect -8309 -3134 -8308 -3114
rect -8306 -3134 -8305 -3114
rect -8257 -3134 -8256 -3114
rect -8254 -3134 -8253 -3114
rect -8205 -3134 -8204 -3114
rect -8202 -3134 -8201 -3114
rect -8153 -3134 -8152 -3114
rect -8150 -3134 -8149 -3114
rect -7870 -3125 -7860 -3124
rect -7766 -3121 -7765 -3111
rect -7763 -3121 -7762 -3111
rect -7730 -3113 -7729 -3103
rect -7727 -3113 -7726 -3103
rect -7870 -3128 -7860 -3127
rect -7607 -3201 -7606 -3181
rect -7604 -3201 -7603 -3181
rect -7564 -3235 -7563 -3224
rect -7561 -3235 -7560 -3224
rect -7607 -3256 -7606 -3236
rect -7604 -3256 -7603 -3236
rect -7462 -3239 -7461 -3219
rect -7459 -3239 -7458 -3219
rect -7269 -3255 -7268 -3235
rect -7266 -3255 -7265 -3235
rect -7419 -3273 -7418 -3262
rect -7416 -3273 -7415 -3262
rect -7462 -3294 -7461 -3274
rect -7459 -3294 -7458 -3274
rect -7123 -3253 -7122 -3233
rect -7120 -3253 -7119 -3233
rect -6979 -3257 -6978 -3237
rect -6976 -3257 -6975 -3237
rect -7226 -3289 -7225 -3278
rect -7223 -3289 -7222 -3278
rect -7080 -3287 -7079 -3276
rect -7077 -3287 -7076 -3276
rect -6824 -3259 -6823 -3239
rect -6821 -3259 -6820 -3239
rect -7269 -3310 -7268 -3290
rect -7266 -3310 -7265 -3290
rect -7123 -3308 -7122 -3288
rect -7120 -3308 -7119 -3288
rect -6936 -3291 -6935 -3280
rect -6933 -3291 -6932 -3280
rect -6689 -3267 -6688 -3247
rect -6686 -3267 -6685 -3247
rect -6979 -3312 -6978 -3292
rect -6976 -3312 -6975 -3292
rect -6781 -3293 -6780 -3282
rect -6778 -3293 -6777 -3282
rect -6824 -3314 -6823 -3294
rect -6821 -3314 -6820 -3294
rect -6646 -3301 -6645 -3290
rect -6643 -3301 -6642 -3290
rect -8094 -3367 -8093 -3347
rect -8091 -3367 -8090 -3347
rect -8062 -3367 -8061 -3347
rect -8059 -3367 -8058 -3347
rect -7825 -3362 -7824 -3342
rect -7822 -3362 -7821 -3342
rect -6689 -3322 -6688 -3302
rect -6686 -3322 -6685 -3302
rect -6498 -3308 -6497 -3298
rect -6495 -3308 -6494 -3298
rect -6562 -3318 -6561 -3308
rect -6559 -3318 -6558 -3308
rect -6529 -3318 -6528 -3308
rect -6526 -3318 -6525 -3308
rect -8191 -3391 -8190 -3371
rect -8188 -3391 -8187 -3371
rect -8139 -3391 -8138 -3371
rect -8136 -3391 -8135 -3371
rect -6336 -3364 -6335 -3354
rect -6333 -3364 -6332 -3354
rect -6400 -3374 -6399 -3364
rect -6397 -3374 -6396 -3364
rect -6367 -3374 -6366 -3364
rect -6364 -3374 -6363 -3364
rect -7782 -3396 -7781 -3385
rect -7779 -3396 -7778 -3385
rect -7825 -3417 -7824 -3397
rect -7822 -3417 -7821 -3397
rect -8295 -3438 -8294 -3418
rect -8292 -3438 -8291 -3418
rect -8243 -3438 -8242 -3418
rect -8240 -3438 -8239 -3418
rect -8191 -3438 -8190 -3418
rect -8188 -3438 -8187 -3418
rect -8139 -3438 -8138 -3418
rect -8136 -3438 -8135 -3418
rect -6178 -3420 -6177 -3410
rect -6175 -3420 -6174 -3410
rect -6242 -3430 -6241 -3420
rect -6239 -3430 -6238 -3420
rect -6209 -3430 -6208 -3420
rect -6206 -3430 -6205 -3420
rect -6012 -3496 -6011 -3486
rect -6009 -3496 -6008 -3486
rect -6076 -3506 -6075 -3496
rect -6073 -3506 -6072 -3496
rect -6043 -3506 -6042 -3496
rect -6040 -3506 -6039 -3496
rect -5708 -3517 -5707 -3497
rect -5705 -3517 -5704 -3497
rect -5676 -3517 -5675 -3497
rect -5673 -3517 -5672 -3497
rect -5805 -3541 -5804 -3521
rect -5802 -3541 -5801 -3521
rect -5753 -3541 -5752 -3521
rect -5750 -3541 -5749 -3521
rect -5541 -3556 -5540 -3545
rect -5538 -3556 -5537 -3545
rect -5909 -3588 -5908 -3568
rect -5906 -3588 -5905 -3568
rect -5857 -3588 -5856 -3568
rect -5854 -3588 -5853 -3568
rect -5805 -3588 -5804 -3568
rect -5802 -3588 -5801 -3568
rect -5753 -3588 -5752 -3568
rect -5750 -3588 -5749 -3568
rect -7864 -3925 -7854 -3924
rect -7864 -3928 -7854 -3927
rect -7760 -3939 -7759 -3931
rect -7757 -3939 -7756 -3931
rect -8039 -3975 -8038 -3955
rect -8036 -3975 -8035 -3955
rect -8007 -3975 -8006 -3955
rect -8004 -3975 -8003 -3955
rect -7864 -3976 -7854 -3975
rect -7760 -3972 -7759 -3962
rect -7757 -3972 -7756 -3962
rect -7724 -3964 -7723 -3954
rect -7721 -3964 -7720 -3954
rect -7864 -3979 -7854 -3978
rect -8136 -3999 -8135 -3979
rect -8133 -3999 -8132 -3979
rect -8084 -3999 -8083 -3979
rect -8081 -3999 -8080 -3979
rect -7599 -4016 -7598 -3996
rect -7596 -4016 -7595 -3996
rect -8240 -4046 -8239 -4026
rect -8237 -4046 -8236 -4026
rect -8188 -4046 -8187 -4026
rect -8185 -4046 -8184 -4026
rect -8136 -4046 -8135 -4026
rect -8133 -4046 -8132 -4026
rect -8084 -4046 -8083 -4026
rect -8081 -4046 -8080 -4026
rect -7430 -4015 -7429 -3995
rect -7427 -4015 -7426 -3995
rect -7266 -4013 -7265 -3993
rect -7263 -4013 -7262 -3993
rect -7126 -4015 -7125 -3995
rect -7123 -4015 -7122 -3995
rect -7556 -4050 -7555 -4039
rect -7553 -4050 -7552 -4039
rect -7387 -4049 -7386 -4038
rect -7384 -4049 -7383 -4038
rect -7223 -4047 -7222 -4036
rect -7220 -4047 -7219 -4036
rect -6975 -4028 -6974 -4008
rect -6972 -4028 -6971 -4008
rect -7599 -4071 -7598 -4051
rect -7596 -4071 -7595 -4051
rect -7430 -4070 -7429 -4050
rect -7427 -4070 -7426 -4050
rect -7266 -4068 -7265 -4048
rect -7263 -4068 -7262 -4048
rect -7083 -4049 -7082 -4038
rect -7080 -4049 -7079 -4038
rect -7126 -4070 -7125 -4050
rect -7123 -4070 -7122 -4050
rect -6932 -4062 -6931 -4051
rect -6929 -4062 -6928 -4051
rect -6635 -4055 -6634 -4045
rect -6632 -4055 -6631 -4045
rect -6975 -4083 -6974 -4063
rect -6972 -4083 -6971 -4063
rect -6699 -4065 -6698 -4055
rect -6696 -4065 -6695 -4055
rect -6666 -4065 -6665 -4055
rect -6663 -4065 -6662 -4055
rect -8022 -4216 -8021 -4196
rect -8019 -4216 -8018 -4196
rect -7990 -4216 -7989 -4196
rect -7987 -4216 -7986 -4196
rect -8119 -4240 -8118 -4220
rect -8116 -4240 -8115 -4220
rect -8067 -4240 -8066 -4220
rect -8064 -4240 -8063 -4220
rect -6812 -4232 -6811 -4212
rect -6809 -4232 -6808 -4212
rect -8223 -4287 -8222 -4267
rect -8220 -4287 -8219 -4267
rect -8171 -4287 -8170 -4267
rect -8168 -4287 -8167 -4267
rect -8119 -4287 -8118 -4267
rect -8116 -4287 -8115 -4267
rect -8067 -4287 -8066 -4267
rect -8064 -4287 -8063 -4267
rect -7832 -4277 -7831 -4257
rect -7829 -4277 -7828 -4257
rect -6769 -4266 -6768 -4255
rect -6766 -4266 -6765 -4255
rect -6501 -4265 -6500 -4255
rect -6498 -4265 -6497 -4255
rect -6812 -4287 -6811 -4267
rect -6809 -4287 -6808 -4267
rect -6565 -4275 -6564 -4265
rect -6562 -4275 -6561 -4265
rect -6532 -4275 -6531 -4265
rect -6529 -4275 -6528 -4265
rect -7789 -4311 -7788 -4300
rect -7786 -4311 -7785 -4300
rect -7832 -4332 -7831 -4312
rect -7829 -4332 -7828 -4312
rect -6197 -4385 -6192 -4379
rect -6193 -4389 -6192 -4385
rect -6190 -4383 -6189 -4379
rect -6190 -4389 -6185 -4383
rect -6354 -4425 -6353 -4415
rect -6351 -4425 -6350 -4415
rect -6418 -4435 -6417 -4425
rect -6415 -4435 -6414 -4425
rect -6385 -4435 -6384 -4425
rect -6382 -4435 -6381 -4425
rect -6197 -4439 -6192 -4433
rect -6193 -4443 -6192 -4439
rect -6190 -4437 -6189 -4433
rect -6190 -4443 -6185 -4437
rect -6175 -4437 -6174 -4433
rect -6179 -4443 -6174 -4437
rect -6172 -4437 -6171 -4433
rect -6172 -4443 -6167 -4437
rect -5875 -4442 -5874 -4422
rect -5872 -4442 -5871 -4422
rect -5843 -4442 -5842 -4422
rect -5840 -4442 -5839 -4422
rect -5972 -4466 -5971 -4446
rect -5969 -4466 -5968 -4446
rect -5920 -4466 -5919 -4446
rect -5917 -4466 -5916 -4446
rect -5717 -4468 -5716 -4457
rect -5714 -4468 -5713 -4457
rect -6076 -4513 -6075 -4493
rect -6073 -4513 -6072 -4493
rect -6024 -4513 -6023 -4493
rect -6021 -4513 -6020 -4493
rect -5972 -4513 -5971 -4493
rect -5969 -4513 -5968 -4493
rect -5920 -4513 -5919 -4493
rect -5917 -4513 -5916 -4493
rect -7864 -4693 -7854 -4692
rect -7864 -4696 -7854 -4695
rect -7760 -4707 -7759 -4699
rect -7757 -4707 -7756 -4699
rect -7864 -4744 -7854 -4743
rect -7760 -4740 -7759 -4730
rect -7757 -4740 -7756 -4730
rect -7724 -4732 -7723 -4722
rect -7721 -4732 -7720 -4722
rect -7864 -4747 -7854 -4746
rect -8033 -4779 -8032 -4759
rect -8030 -4779 -8029 -4759
rect -8001 -4779 -8000 -4759
rect -7998 -4779 -7997 -4759
rect -8130 -4803 -8129 -4783
rect -8127 -4803 -8126 -4783
rect -8078 -4803 -8077 -4783
rect -8075 -4803 -8074 -4783
rect -7578 -4789 -7577 -4769
rect -7575 -4789 -7574 -4769
rect -7535 -4823 -7534 -4812
rect -7532 -4823 -7531 -4812
rect -8234 -4850 -8233 -4830
rect -8231 -4850 -8230 -4830
rect -8182 -4850 -8181 -4830
rect -8179 -4850 -8178 -4830
rect -8130 -4850 -8129 -4830
rect -8127 -4850 -8126 -4830
rect -8078 -4850 -8077 -4830
rect -8075 -4850 -8074 -4830
rect -7578 -4844 -7577 -4824
rect -7575 -4844 -7574 -4824
rect -7382 -4915 -7381 -4905
rect -7379 -4915 -7378 -4905
rect -7446 -4925 -7445 -4915
rect -7443 -4925 -7442 -4915
rect -7413 -4925 -7412 -4915
rect -7410 -4925 -7409 -4915
rect -7577 -4994 -7576 -4974
rect -7574 -4994 -7573 -4974
rect -7534 -5028 -7533 -5017
rect -7531 -5028 -7530 -5017
rect -7115 -4996 -7110 -4990
rect -7111 -5000 -7110 -4996
rect -7108 -4994 -7107 -4990
rect -7108 -5000 -7103 -4994
rect -7236 -5028 -7235 -5018
rect -7233 -5028 -7232 -5018
rect -7577 -5049 -7576 -5029
rect -7574 -5049 -7573 -5029
rect -7300 -5038 -7299 -5028
rect -7297 -5038 -7296 -5028
rect -7267 -5038 -7266 -5028
rect -7264 -5038 -7263 -5028
rect -7115 -5050 -7110 -5044
rect -8020 -5091 -8019 -5071
rect -8017 -5091 -8016 -5071
rect -7988 -5091 -7987 -5071
rect -7985 -5091 -7984 -5071
rect -7111 -5054 -7110 -5050
rect -7108 -5048 -7107 -5044
rect -7108 -5054 -7103 -5048
rect -7093 -5048 -7092 -5044
rect -7097 -5054 -7092 -5048
rect -7090 -5048 -7089 -5044
rect -7090 -5054 -7085 -5048
rect -8117 -5115 -8116 -5095
rect -8114 -5115 -8113 -5095
rect -8065 -5115 -8064 -5095
rect -8062 -5115 -8061 -5095
rect -6794 -5051 -6793 -5031
rect -6791 -5051 -6790 -5031
rect -6762 -5051 -6761 -5031
rect -6759 -5051 -6758 -5031
rect -6891 -5075 -6890 -5055
rect -6888 -5075 -6887 -5055
rect -6839 -5075 -6838 -5055
rect -6836 -5075 -6835 -5055
rect -7838 -5126 -7837 -5106
rect -7835 -5126 -7834 -5106
rect -6683 -5088 -6682 -5077
rect -6680 -5088 -6679 -5077
rect -3990 -5096 -3985 -5090
rect -3986 -5100 -3985 -5096
rect -3983 -5094 -3982 -5090
rect -3983 -5100 -3978 -5094
rect -6995 -5122 -6994 -5102
rect -6992 -5122 -6991 -5102
rect -6943 -5122 -6942 -5102
rect -6940 -5122 -6939 -5102
rect -6891 -5122 -6890 -5102
rect -6888 -5122 -6887 -5102
rect -6839 -5122 -6838 -5102
rect -6836 -5122 -6835 -5102
rect -8221 -5162 -8220 -5142
rect -8218 -5162 -8217 -5142
rect -8169 -5162 -8168 -5142
rect -8166 -5162 -8165 -5142
rect -8117 -5162 -8116 -5142
rect -8114 -5162 -8113 -5142
rect -8065 -5162 -8064 -5142
rect -8062 -5162 -8061 -5142
rect -7795 -5160 -7794 -5149
rect -7792 -5160 -7791 -5149
rect -3990 -5150 -3985 -5144
rect -3986 -5154 -3985 -5150
rect -3983 -5148 -3982 -5144
rect -3983 -5154 -3978 -5148
rect -3968 -5148 -3967 -5144
rect -3972 -5154 -3967 -5148
rect -3965 -5148 -3964 -5144
rect -3965 -5154 -3960 -5148
rect -7838 -5181 -7837 -5161
rect -7835 -5181 -7834 -5161
rect -7886 -5455 -7876 -5454
rect -7886 -5458 -7876 -5457
rect -8033 -5485 -8032 -5465
rect -8030 -5485 -8029 -5465
rect -8001 -5485 -8000 -5465
rect -7998 -5485 -7997 -5465
rect -7782 -5469 -7781 -5461
rect -7779 -5469 -7778 -5461
rect -8130 -5509 -8129 -5489
rect -8127 -5509 -8126 -5489
rect -8078 -5509 -8077 -5489
rect -8075 -5509 -8074 -5489
rect -7886 -5506 -7876 -5505
rect -7782 -5502 -7781 -5492
rect -7779 -5502 -7778 -5492
rect -7746 -5494 -7745 -5484
rect -7743 -5494 -7742 -5484
rect -7886 -5509 -7876 -5508
rect -8234 -5556 -8233 -5536
rect -8231 -5556 -8230 -5536
rect -8182 -5556 -8181 -5536
rect -8179 -5556 -8178 -5536
rect -8130 -5556 -8129 -5536
rect -8127 -5556 -8126 -5536
rect -8078 -5556 -8077 -5536
rect -8075 -5556 -8074 -5536
rect -7666 -5569 -7665 -5549
rect -7663 -5569 -7662 -5549
rect -7623 -5603 -7622 -5592
rect -7620 -5603 -7619 -5592
rect -7666 -5624 -7665 -5604
rect -7663 -5624 -7662 -5604
rect -8030 -5734 -8029 -5714
rect -8027 -5734 -8026 -5714
rect -7998 -5734 -7997 -5714
rect -7995 -5734 -7994 -5714
rect -8127 -5758 -8126 -5738
rect -8124 -5758 -8123 -5738
rect -8075 -5758 -8074 -5738
rect -8072 -5758 -8071 -5738
rect -7835 -5749 -7834 -5729
rect -7832 -5749 -7831 -5729
rect -7307 -5720 -7302 -5714
rect -7303 -5724 -7302 -5720
rect -7300 -5718 -7299 -5714
rect -7300 -5724 -7295 -5718
rect -6978 -5705 -6977 -5685
rect -6975 -5705 -6974 -5685
rect -6946 -5705 -6945 -5685
rect -6943 -5705 -6942 -5685
rect -7075 -5729 -7074 -5709
rect -7072 -5729 -7071 -5709
rect -7023 -5729 -7022 -5709
rect -7020 -5729 -7019 -5709
rect -7488 -5758 -7487 -5748
rect -7485 -5758 -7484 -5748
rect -7552 -5768 -7551 -5758
rect -7549 -5768 -7548 -5758
rect -7519 -5768 -7518 -5758
rect -7516 -5768 -7515 -5758
rect -7792 -5783 -7791 -5772
rect -7789 -5783 -7788 -5772
rect -7307 -5774 -7302 -5768
rect -7303 -5778 -7302 -5774
rect -7300 -5772 -7299 -5768
rect -7300 -5778 -7295 -5772
rect -7285 -5772 -7284 -5768
rect -7289 -5778 -7284 -5772
rect -7282 -5772 -7281 -5768
rect -7282 -5778 -7277 -5772
rect -7179 -5776 -7178 -5756
rect -7176 -5776 -7175 -5756
rect -7127 -5776 -7126 -5756
rect -7124 -5776 -7123 -5756
rect -7075 -5776 -7074 -5756
rect -7072 -5776 -7071 -5756
rect -7023 -5776 -7022 -5756
rect -7020 -5776 -7019 -5756
rect -6819 -5763 -6818 -5752
rect -6816 -5763 -6815 -5752
rect -8231 -5805 -8230 -5785
rect -8228 -5805 -8227 -5785
rect -8179 -5805 -8178 -5785
rect -8176 -5805 -8175 -5785
rect -8127 -5805 -8126 -5785
rect -8124 -5805 -8123 -5785
rect -8075 -5805 -8074 -5785
rect -8072 -5805 -8071 -5785
rect -7835 -5804 -7834 -5784
rect -7832 -5804 -7831 -5784
rect -7635 -5836 -7630 -5830
rect -7631 -5840 -7630 -5836
rect -7628 -5834 -7627 -5830
rect -7628 -5840 -7623 -5834
rect -7635 -5890 -7630 -5884
rect -7631 -5894 -7630 -5890
rect -7628 -5888 -7627 -5884
rect -7628 -5894 -7623 -5888
rect -7613 -5888 -7612 -5884
rect -7617 -5894 -7612 -5888
rect -7610 -5888 -7609 -5884
rect -7610 -5894 -7605 -5888
rect -7255 -5945 -7254 -5925
rect -7252 -5945 -7251 -5925
rect -7223 -5945 -7222 -5925
rect -7220 -5945 -7219 -5925
rect -7352 -5969 -7351 -5949
rect -7349 -5969 -7348 -5949
rect -7300 -5969 -7299 -5949
rect -7297 -5969 -7296 -5949
rect -7120 -5985 -7119 -5974
rect -7117 -5985 -7116 -5974
rect -7456 -6016 -7455 -5996
rect -7453 -6016 -7452 -5996
rect -7404 -6016 -7403 -5996
rect -7401 -6016 -7400 -5996
rect -7352 -6016 -7351 -5996
rect -7349 -6016 -7348 -5996
rect -7300 -6016 -7299 -5996
rect -7297 -6016 -7296 -5996
rect -7655 -6045 -7654 -6025
rect -7652 -6045 -7651 -6025
rect -7623 -6045 -7622 -6025
rect -7620 -6045 -7619 -6025
rect -7752 -6069 -7751 -6049
rect -7749 -6069 -7748 -6049
rect -7700 -6069 -7699 -6049
rect -7697 -6069 -7696 -6049
rect -7856 -6116 -7855 -6096
rect -7853 -6116 -7852 -6096
rect -7804 -6116 -7803 -6096
rect -7801 -6116 -7800 -6096
rect -7752 -6116 -7751 -6096
rect -7749 -6116 -7748 -6096
rect -7700 -6116 -7699 -6096
rect -7697 -6116 -7696 -6096
rect -7544 -6230 -7543 -6219
rect -7541 -6230 -7540 -6219
<< pdiffusion >>
rect -2914 -530 -2913 -510
rect -2911 -530 -2910 -510
rect -2887 -530 -2886 -510
rect -2884 -530 -2883 -510
rect -2852 -600 -2851 -560
rect -2849 -600 -2848 -560
rect -2540 -601 -2520 -600
rect -2540 -604 -2520 -603
rect -2438 -612 -2437 -592
rect -2435 -612 -2434 -592
rect -2540 -652 -2520 -651
rect -2540 -655 -2520 -654
rect -2284 -678 -2283 -658
rect -2281 -678 -2280 -658
rect -2284 -725 -2283 -706
rect -2281 -725 -2280 -706
rect -2235 -722 -2234 -702
rect -2232 -722 -2231 -702
rect -1986 -708 -1985 -668
rect -1983 -708 -1982 -668
rect -1934 -708 -1933 -668
rect -1931 -708 -1930 -668
rect -1882 -708 -1881 -668
rect -1879 -708 -1878 -668
rect -1830 -708 -1829 -668
rect -1827 -708 -1826 -668
rect -1785 -700 -1784 -660
rect -1782 -700 -1781 -660
rect -1753 -700 -1752 -660
rect -1750 -700 -1749 -660
rect -1986 -770 -1985 -730
rect -1983 -770 -1982 -730
rect -1934 -770 -1933 -730
rect -1931 -770 -1930 -730
rect -8309 -3031 -8308 -2991
rect -8306 -3031 -8305 -2991
rect -8257 -3031 -8256 -2991
rect -8254 -3031 -8253 -2991
rect -8205 -3031 -8204 -2991
rect -8202 -3031 -8201 -2991
rect -8153 -3031 -8152 -2991
rect -8150 -3031 -8149 -2991
rect -8108 -3023 -8107 -2983
rect -8105 -3023 -8104 -2983
rect -8076 -3023 -8075 -2983
rect -8073 -3023 -8072 -2983
rect -8309 -3093 -8308 -3053
rect -8306 -3093 -8305 -3053
rect -8257 -3093 -8256 -3053
rect -8254 -3093 -8253 -3053
rect -7832 -3074 -7812 -3073
rect -7832 -3077 -7812 -3076
rect -7730 -3085 -7729 -3065
rect -7727 -3085 -7726 -3065
rect -7832 -3125 -7812 -3124
rect -7832 -3128 -7812 -3127
rect -7626 -3127 -7625 -3107
rect -7623 -3127 -7622 -3107
rect -7599 -3127 -7598 -3107
rect -7596 -3127 -7595 -3107
rect -7564 -3197 -7563 -3157
rect -7561 -3197 -7560 -3157
rect -7481 -3165 -7480 -3145
rect -7478 -3165 -7477 -3145
rect -7454 -3165 -7453 -3145
rect -7451 -3165 -7450 -3145
rect -7288 -3181 -7287 -3161
rect -7285 -3181 -7284 -3161
rect -7261 -3181 -7260 -3161
rect -7258 -3181 -7257 -3161
rect -7142 -3179 -7141 -3159
rect -7139 -3179 -7138 -3159
rect -7115 -3179 -7114 -3159
rect -7112 -3179 -7111 -3159
rect -7419 -3235 -7418 -3195
rect -7416 -3235 -7415 -3195
rect -6998 -3183 -6997 -3163
rect -6995 -3183 -6994 -3163
rect -6971 -3183 -6970 -3163
rect -6968 -3183 -6967 -3163
rect -7226 -3251 -7225 -3211
rect -7223 -3251 -7222 -3211
rect -6843 -3185 -6842 -3165
rect -6840 -3185 -6839 -3165
rect -6816 -3185 -6815 -3165
rect -6813 -3185 -6812 -3165
rect -8295 -3335 -8294 -3295
rect -8292 -3335 -8291 -3295
rect -8243 -3335 -8242 -3295
rect -8240 -3335 -8239 -3295
rect -8191 -3335 -8190 -3295
rect -8188 -3335 -8187 -3295
rect -8139 -3335 -8138 -3295
rect -8136 -3335 -8135 -3295
rect -8094 -3327 -8093 -3287
rect -8091 -3327 -8090 -3287
rect -8062 -3327 -8061 -3287
rect -8059 -3327 -8058 -3287
rect -7844 -3288 -7843 -3268
rect -7841 -3288 -7840 -3268
rect -7817 -3288 -7816 -3268
rect -7814 -3288 -7813 -3268
rect -7080 -3249 -7079 -3209
rect -7077 -3249 -7076 -3209
rect -6708 -3193 -6707 -3173
rect -6705 -3193 -6704 -3173
rect -6681 -3193 -6680 -3173
rect -6678 -3193 -6677 -3173
rect -6936 -3253 -6935 -3213
rect -6933 -3253 -6932 -3213
rect -6781 -3255 -6780 -3215
rect -6778 -3255 -6777 -3215
rect -6646 -3263 -6645 -3223
rect -6643 -3263 -6642 -3223
rect -6547 -3236 -6546 -3216
rect -6544 -3236 -6543 -3216
rect -6547 -3283 -6546 -3264
rect -6544 -3283 -6543 -3264
rect -8295 -3397 -8294 -3357
rect -8292 -3397 -8291 -3357
rect -8243 -3397 -8242 -3357
rect -8240 -3397 -8239 -3357
rect -7782 -3358 -7781 -3318
rect -7779 -3358 -7778 -3318
rect -6498 -3280 -6497 -3260
rect -6495 -3280 -6494 -3260
rect -6385 -3292 -6384 -3272
rect -6382 -3292 -6381 -3272
rect -6385 -3339 -6384 -3320
rect -6382 -3339 -6381 -3320
rect -6336 -3336 -6335 -3316
rect -6333 -3336 -6332 -3316
rect -6227 -3348 -6226 -3328
rect -6224 -3348 -6223 -3328
rect -6227 -3395 -6226 -3376
rect -6224 -3395 -6223 -3376
rect -6178 -3392 -6177 -3372
rect -6175 -3392 -6174 -3372
rect -6061 -3424 -6060 -3404
rect -6058 -3424 -6057 -3404
rect -6061 -3471 -6060 -3452
rect -6058 -3471 -6057 -3452
rect -6012 -3468 -6011 -3448
rect -6009 -3468 -6008 -3448
rect -5909 -3485 -5908 -3445
rect -5906 -3485 -5905 -3445
rect -5857 -3485 -5856 -3445
rect -5854 -3485 -5853 -3445
rect -5805 -3485 -5804 -3445
rect -5802 -3485 -5801 -3445
rect -5753 -3485 -5752 -3445
rect -5750 -3485 -5749 -3445
rect -5708 -3477 -5707 -3437
rect -5705 -3477 -5704 -3437
rect -5676 -3477 -5675 -3437
rect -5673 -3477 -5672 -3437
rect -5909 -3547 -5908 -3507
rect -5906 -3547 -5905 -3507
rect -5857 -3547 -5856 -3507
rect -5854 -3547 -5853 -3507
rect -5541 -3518 -5540 -3478
rect -5538 -3518 -5537 -3478
rect -8240 -3943 -8239 -3903
rect -8237 -3943 -8236 -3903
rect -8188 -3943 -8187 -3903
rect -8185 -3943 -8184 -3903
rect -8136 -3943 -8135 -3903
rect -8133 -3943 -8132 -3903
rect -8084 -3943 -8083 -3903
rect -8081 -3943 -8080 -3903
rect -8039 -3935 -8038 -3895
rect -8036 -3935 -8035 -3895
rect -8007 -3935 -8006 -3895
rect -8004 -3935 -8003 -3895
rect -7826 -3925 -7806 -3924
rect -7826 -3928 -7806 -3927
rect -7724 -3936 -7723 -3916
rect -7721 -3936 -7720 -3916
rect -8240 -4005 -8239 -3965
rect -8237 -4005 -8236 -3965
rect -8188 -4005 -8187 -3965
rect -8185 -4005 -8184 -3965
rect -7618 -3942 -7617 -3922
rect -7615 -3942 -7614 -3922
rect -7591 -3942 -7590 -3922
rect -7588 -3942 -7587 -3922
rect -7449 -3941 -7448 -3921
rect -7446 -3941 -7445 -3921
rect -7422 -3941 -7421 -3921
rect -7419 -3941 -7418 -3921
rect -7285 -3939 -7284 -3919
rect -7282 -3939 -7281 -3919
rect -7258 -3939 -7257 -3919
rect -7255 -3939 -7254 -3919
rect -7145 -3941 -7144 -3921
rect -7142 -3941 -7141 -3921
rect -7118 -3941 -7117 -3921
rect -7115 -3941 -7114 -3921
rect -6994 -3954 -6993 -3934
rect -6991 -3954 -6990 -3934
rect -6967 -3954 -6966 -3934
rect -6964 -3954 -6963 -3934
rect -7826 -3976 -7806 -3975
rect -7826 -3979 -7806 -3978
rect -7556 -4012 -7555 -3972
rect -7553 -4012 -7552 -3972
rect -7387 -4011 -7386 -3971
rect -7384 -4011 -7383 -3971
rect -7223 -4009 -7222 -3969
rect -7220 -4009 -7219 -3969
rect -7083 -4011 -7082 -3971
rect -7080 -4011 -7079 -3971
rect -6684 -3983 -6683 -3963
rect -6681 -3983 -6680 -3963
rect -6932 -4024 -6931 -3984
rect -6929 -4024 -6928 -3984
rect -6684 -4030 -6683 -4011
rect -6681 -4030 -6680 -4011
rect -6635 -4027 -6634 -4007
rect -6632 -4027 -6631 -4007
rect -8223 -4184 -8222 -4144
rect -8220 -4184 -8219 -4144
rect -8171 -4184 -8170 -4144
rect -8168 -4184 -8167 -4144
rect -8119 -4184 -8118 -4144
rect -8116 -4184 -8115 -4144
rect -8067 -4184 -8066 -4144
rect -8064 -4184 -8063 -4144
rect -8022 -4176 -8021 -4136
rect -8019 -4176 -8018 -4136
rect -7990 -4176 -7989 -4136
rect -7987 -4176 -7986 -4136
rect -6831 -4158 -6830 -4138
rect -6828 -4158 -6827 -4138
rect -6804 -4158 -6803 -4138
rect -6801 -4158 -6800 -4138
rect -8223 -4246 -8222 -4206
rect -8220 -4246 -8219 -4206
rect -8171 -4246 -8170 -4206
rect -8168 -4246 -8167 -4206
rect -7851 -4203 -7850 -4183
rect -7848 -4203 -7847 -4183
rect -7824 -4203 -7823 -4183
rect -7821 -4203 -7820 -4183
rect -6769 -4228 -6768 -4188
rect -6766 -4228 -6765 -4188
rect -6550 -4193 -6549 -4173
rect -6547 -4193 -6546 -4173
rect -7789 -4273 -7788 -4233
rect -7786 -4273 -7785 -4233
rect -6550 -4240 -6549 -4221
rect -6547 -4240 -6546 -4221
rect -6501 -4237 -6500 -4217
rect -6498 -4237 -6497 -4217
rect -6403 -4353 -6402 -4333
rect -6400 -4353 -6399 -4333
rect -6193 -4350 -6192 -4346
rect -6403 -4400 -6402 -4381
rect -6400 -4400 -6399 -4381
rect -6197 -4366 -6192 -4350
rect -6190 -4362 -6185 -4346
rect -6190 -4366 -6189 -4362
rect -6354 -4397 -6353 -4377
rect -6351 -4397 -6350 -4377
rect -6193 -4405 -6192 -4401
rect -6197 -4421 -6192 -4405
rect -6190 -4417 -6185 -4401
rect -6190 -4421 -6189 -4417
rect -6179 -4417 -6174 -4401
rect -6175 -4421 -6174 -4417
rect -6172 -4417 -6167 -4401
rect -6076 -4410 -6075 -4370
rect -6073 -4410 -6072 -4370
rect -6024 -4410 -6023 -4370
rect -6021 -4410 -6020 -4370
rect -5972 -4410 -5971 -4370
rect -5969 -4410 -5968 -4370
rect -5920 -4410 -5919 -4370
rect -5917 -4410 -5916 -4370
rect -5875 -4402 -5874 -4362
rect -5872 -4402 -5871 -4362
rect -5843 -4402 -5842 -4362
rect -5840 -4402 -5839 -4362
rect -6172 -4421 -6171 -4417
rect -6076 -4472 -6075 -4432
rect -6073 -4472 -6072 -4432
rect -6024 -4472 -6023 -4432
rect -6021 -4472 -6020 -4432
rect -5717 -4430 -5716 -4390
rect -5714 -4430 -5713 -4390
rect -7826 -4693 -7806 -4692
rect -8234 -4747 -8233 -4707
rect -8231 -4747 -8230 -4707
rect -8182 -4747 -8181 -4707
rect -8179 -4747 -8178 -4707
rect -8130 -4747 -8129 -4707
rect -8127 -4747 -8126 -4707
rect -8078 -4747 -8077 -4707
rect -8075 -4747 -8074 -4707
rect -8033 -4739 -8032 -4699
rect -8030 -4739 -8029 -4699
rect -8001 -4739 -8000 -4699
rect -7998 -4739 -7997 -4699
rect -7826 -4696 -7806 -4695
rect -7724 -4704 -7723 -4684
rect -7721 -4704 -7720 -4684
rect -7597 -4715 -7596 -4695
rect -7594 -4715 -7593 -4695
rect -7570 -4715 -7569 -4695
rect -7567 -4715 -7566 -4695
rect -7826 -4744 -7806 -4743
rect -7826 -4747 -7806 -4746
rect -8234 -4809 -8233 -4769
rect -8231 -4809 -8230 -4769
rect -8182 -4809 -8181 -4769
rect -8179 -4809 -8178 -4769
rect -7535 -4785 -7534 -4745
rect -7532 -4785 -7531 -4745
rect -7431 -4843 -7430 -4823
rect -7428 -4843 -7427 -4823
rect -7431 -4890 -7430 -4871
rect -7428 -4890 -7427 -4871
rect -7596 -4920 -7595 -4900
rect -7593 -4920 -7592 -4900
rect -7569 -4920 -7568 -4900
rect -7566 -4920 -7565 -4900
rect -7382 -4887 -7381 -4867
rect -7379 -4887 -7378 -4867
rect -7534 -4990 -7533 -4950
rect -7531 -4990 -7530 -4950
rect -7285 -4956 -7284 -4936
rect -7282 -4956 -7281 -4936
rect -7111 -4961 -7110 -4957
rect -8221 -5059 -8220 -5019
rect -8218 -5059 -8217 -5019
rect -8169 -5059 -8168 -5019
rect -8166 -5059 -8165 -5019
rect -8117 -5059 -8116 -5019
rect -8114 -5059 -8113 -5019
rect -8065 -5059 -8064 -5019
rect -8062 -5059 -8061 -5019
rect -8020 -5051 -8019 -5011
rect -8017 -5051 -8016 -5011
rect -7988 -5051 -7987 -5011
rect -7985 -5051 -7984 -5011
rect -7285 -5003 -7284 -4984
rect -7282 -5003 -7281 -4984
rect -7115 -4977 -7110 -4961
rect -7108 -4973 -7103 -4957
rect -7108 -4977 -7107 -4973
rect -7236 -5000 -7235 -4980
rect -7233 -5000 -7232 -4980
rect -7111 -5016 -7110 -5012
rect -7857 -5052 -7856 -5032
rect -7854 -5052 -7853 -5032
rect -7830 -5052 -7829 -5032
rect -7827 -5052 -7826 -5032
rect -7115 -5032 -7110 -5016
rect -7108 -5028 -7103 -5012
rect -7108 -5032 -7107 -5028
rect -7097 -5028 -7092 -5012
rect -7093 -5032 -7092 -5028
rect -7090 -5028 -7085 -5012
rect -6995 -5019 -6994 -4979
rect -6992 -5019 -6991 -4979
rect -6943 -5019 -6942 -4979
rect -6940 -5019 -6939 -4979
rect -6891 -5019 -6890 -4979
rect -6888 -5019 -6887 -4979
rect -6839 -5019 -6838 -4979
rect -6836 -5019 -6835 -4979
rect -6794 -5011 -6793 -4971
rect -6791 -5011 -6790 -4971
rect -6762 -5011 -6761 -4971
rect -6759 -5011 -6758 -4971
rect -7090 -5032 -7089 -5028
rect -8221 -5121 -8220 -5081
rect -8218 -5121 -8217 -5081
rect -8169 -5121 -8168 -5081
rect -8166 -5121 -8165 -5081
rect -6995 -5081 -6994 -5041
rect -6992 -5081 -6991 -5041
rect -6943 -5081 -6942 -5041
rect -6940 -5081 -6939 -5041
rect -6683 -5050 -6682 -5010
rect -6680 -5050 -6679 -5010
rect -3986 -5061 -3985 -5057
rect -3990 -5077 -3985 -5061
rect -3983 -5073 -3978 -5057
rect -3983 -5077 -3982 -5073
rect -7795 -5122 -7794 -5082
rect -7792 -5122 -7791 -5082
rect -3986 -5116 -3985 -5112
rect -3990 -5132 -3985 -5116
rect -3983 -5128 -3978 -5112
rect -3983 -5132 -3982 -5128
rect -3972 -5128 -3967 -5112
rect -3968 -5132 -3967 -5128
rect -3965 -5128 -3960 -5112
rect -3965 -5132 -3964 -5128
rect -8234 -5453 -8233 -5413
rect -8231 -5453 -8230 -5413
rect -8182 -5453 -8181 -5413
rect -8179 -5453 -8178 -5413
rect -8130 -5453 -8129 -5413
rect -8127 -5453 -8126 -5413
rect -8078 -5453 -8077 -5413
rect -8075 -5453 -8074 -5413
rect -8033 -5445 -8032 -5405
rect -8030 -5445 -8029 -5405
rect -8001 -5445 -8000 -5405
rect -7998 -5445 -7997 -5405
rect -7848 -5455 -7828 -5454
rect -7848 -5458 -7828 -5457
rect -8234 -5515 -8233 -5475
rect -8231 -5515 -8230 -5475
rect -8182 -5515 -8181 -5475
rect -8179 -5515 -8178 -5475
rect -7746 -5466 -7745 -5446
rect -7743 -5466 -7742 -5446
rect -7685 -5495 -7684 -5475
rect -7682 -5495 -7681 -5475
rect -7658 -5495 -7657 -5475
rect -7655 -5495 -7654 -5475
rect -7848 -5506 -7828 -5505
rect -7848 -5509 -7828 -5508
rect -7623 -5565 -7622 -5525
rect -7620 -5565 -7619 -5525
rect -8231 -5702 -8230 -5662
rect -8228 -5702 -8227 -5662
rect -8179 -5702 -8178 -5662
rect -8176 -5702 -8175 -5662
rect -8127 -5702 -8126 -5662
rect -8124 -5702 -8123 -5662
rect -8075 -5702 -8074 -5662
rect -8072 -5702 -8071 -5662
rect -8030 -5694 -8029 -5654
rect -8027 -5694 -8026 -5654
rect -7998 -5694 -7997 -5654
rect -7995 -5694 -7994 -5654
rect -7854 -5675 -7853 -5655
rect -7851 -5675 -7850 -5655
rect -7827 -5675 -7826 -5655
rect -7824 -5675 -7823 -5655
rect -7537 -5686 -7536 -5666
rect -7534 -5686 -7533 -5666
rect -7179 -5673 -7178 -5633
rect -7176 -5673 -7175 -5633
rect -7127 -5673 -7126 -5633
rect -7124 -5673 -7123 -5633
rect -7075 -5673 -7074 -5633
rect -7072 -5673 -7071 -5633
rect -7023 -5673 -7022 -5633
rect -7020 -5673 -7019 -5633
rect -6978 -5665 -6977 -5625
rect -6975 -5665 -6974 -5625
rect -6946 -5665 -6945 -5625
rect -6943 -5665 -6942 -5625
rect -7303 -5685 -7302 -5681
rect -8231 -5764 -8230 -5724
rect -8228 -5764 -8227 -5724
rect -8179 -5764 -8178 -5724
rect -8176 -5764 -8175 -5724
rect -7792 -5745 -7791 -5705
rect -7789 -5745 -7788 -5705
rect -7537 -5733 -7536 -5714
rect -7534 -5733 -7533 -5714
rect -7307 -5701 -7302 -5685
rect -7300 -5697 -7295 -5681
rect -7300 -5701 -7299 -5697
rect -7488 -5730 -7487 -5710
rect -7485 -5730 -7484 -5710
rect -7179 -5735 -7178 -5695
rect -7176 -5735 -7175 -5695
rect -7127 -5735 -7126 -5695
rect -7124 -5735 -7123 -5695
rect -6819 -5725 -6818 -5685
rect -6816 -5725 -6815 -5685
rect -7303 -5740 -7302 -5736
rect -7307 -5756 -7302 -5740
rect -7300 -5752 -7295 -5736
rect -7300 -5756 -7299 -5752
rect -7289 -5752 -7284 -5736
rect -7285 -5756 -7284 -5752
rect -7282 -5752 -7277 -5736
rect -7282 -5756 -7281 -5752
rect -7631 -5801 -7630 -5797
rect -7635 -5817 -7630 -5801
rect -7628 -5813 -7623 -5797
rect -7628 -5817 -7627 -5813
rect -7631 -5856 -7630 -5852
rect -7635 -5872 -7630 -5856
rect -7628 -5868 -7623 -5852
rect -7628 -5872 -7627 -5868
rect -7617 -5868 -7612 -5852
rect -7613 -5872 -7612 -5868
rect -7610 -5868 -7605 -5852
rect -7610 -5872 -7609 -5868
rect -7456 -5913 -7455 -5873
rect -7453 -5913 -7452 -5873
rect -7404 -5913 -7403 -5873
rect -7401 -5913 -7400 -5873
rect -7352 -5913 -7351 -5873
rect -7349 -5913 -7348 -5873
rect -7300 -5913 -7299 -5873
rect -7297 -5913 -7296 -5873
rect -7255 -5905 -7254 -5865
rect -7252 -5905 -7251 -5865
rect -7223 -5905 -7222 -5865
rect -7220 -5905 -7219 -5865
rect -7856 -6013 -7855 -5973
rect -7853 -6013 -7852 -5973
rect -7804 -6013 -7803 -5973
rect -7801 -6013 -7800 -5973
rect -7752 -6013 -7751 -5973
rect -7749 -6013 -7748 -5973
rect -7700 -6013 -7699 -5973
rect -7697 -6013 -7696 -5973
rect -7655 -6005 -7654 -5965
rect -7652 -6005 -7651 -5965
rect -7623 -6005 -7622 -5965
rect -7620 -6005 -7619 -5965
rect -7456 -5975 -7455 -5935
rect -7453 -5975 -7452 -5935
rect -7404 -5975 -7403 -5935
rect -7401 -5975 -7400 -5935
rect -7120 -5947 -7119 -5907
rect -7117 -5947 -7116 -5907
rect -7856 -6075 -7855 -6035
rect -7853 -6075 -7852 -6035
rect -7804 -6075 -7803 -6035
rect -7801 -6075 -7800 -6035
rect -7544 -6192 -7543 -6152
rect -7541 -6192 -7540 -6152
<< ndcontact >>
rect -2899 -604 -2895 -584
rect -2891 -604 -2887 -584
rect -2578 -600 -2568 -596
rect -2578 -608 -2568 -604
rect -2478 -615 -2474 -605
rect -2470 -615 -2466 -605
rect -2856 -638 -2852 -627
rect -2848 -638 -2844 -627
rect -2899 -659 -2895 -639
rect -2891 -659 -2887 -639
rect -2578 -651 -2568 -647
rect -2478 -648 -2474 -638
rect -2470 -648 -2466 -638
rect -2442 -640 -2438 -630
rect -2434 -640 -2430 -630
rect -2578 -659 -2568 -655
rect -2239 -750 -2235 -740
rect -2231 -750 -2227 -740
rect -2303 -760 -2299 -750
rect -2295 -760 -2291 -750
rect -2270 -760 -2266 -750
rect -2262 -760 -2258 -750
rect -1789 -740 -1785 -720
rect -1781 -740 -1777 -720
rect -1757 -740 -1753 -720
rect -1749 -740 -1745 -720
rect -1886 -764 -1882 -744
rect -1878 -764 -1874 -744
rect -1834 -764 -1830 -744
rect -1826 -764 -1822 -744
rect -1990 -811 -1986 -791
rect -1982 -811 -1978 -791
rect -1938 -811 -1934 -791
rect -1930 -811 -1926 -791
rect -1886 -811 -1882 -791
rect -1878 -811 -1874 -791
rect -1834 -811 -1830 -791
rect -1826 -811 -1822 -791
rect -8112 -3063 -8108 -3043
rect -8104 -3063 -8100 -3043
rect -8080 -3063 -8076 -3043
rect -8072 -3063 -8068 -3043
rect -8209 -3087 -8205 -3067
rect -8201 -3087 -8197 -3067
rect -8157 -3087 -8153 -3067
rect -8149 -3087 -8145 -3067
rect -7870 -3073 -7860 -3069
rect -7870 -3081 -7860 -3077
rect -7770 -3088 -7766 -3080
rect -7762 -3088 -7758 -3080
rect -8313 -3134 -8309 -3114
rect -8305 -3134 -8301 -3114
rect -8261 -3134 -8257 -3114
rect -8253 -3134 -8249 -3114
rect -8209 -3134 -8205 -3114
rect -8201 -3134 -8197 -3114
rect -8157 -3134 -8153 -3114
rect -8149 -3134 -8145 -3114
rect -7870 -3124 -7860 -3120
rect -7770 -3121 -7766 -3111
rect -7762 -3121 -7758 -3111
rect -7734 -3113 -7730 -3103
rect -7726 -3113 -7722 -3103
rect -7870 -3132 -7860 -3128
rect -7611 -3201 -7607 -3181
rect -7603 -3201 -7599 -3181
rect -7568 -3235 -7564 -3224
rect -7560 -3235 -7556 -3224
rect -7611 -3256 -7607 -3236
rect -7603 -3256 -7599 -3236
rect -7466 -3239 -7462 -3219
rect -7458 -3239 -7454 -3219
rect -7273 -3255 -7269 -3235
rect -7265 -3255 -7261 -3235
rect -7423 -3273 -7419 -3262
rect -7415 -3273 -7411 -3262
rect -7466 -3294 -7462 -3274
rect -7458 -3294 -7454 -3274
rect -7127 -3253 -7123 -3233
rect -7119 -3253 -7115 -3233
rect -6983 -3257 -6979 -3237
rect -6975 -3257 -6971 -3237
rect -7230 -3289 -7226 -3278
rect -7222 -3289 -7218 -3278
rect -7084 -3287 -7080 -3276
rect -7076 -3287 -7072 -3276
rect -6828 -3259 -6824 -3239
rect -6820 -3259 -6816 -3239
rect -7273 -3310 -7269 -3290
rect -7265 -3310 -7261 -3290
rect -7127 -3308 -7123 -3288
rect -7119 -3308 -7115 -3288
rect -6940 -3291 -6936 -3280
rect -6932 -3291 -6928 -3280
rect -6693 -3267 -6689 -3247
rect -6685 -3267 -6681 -3247
rect -6983 -3312 -6979 -3292
rect -6975 -3312 -6971 -3292
rect -6785 -3293 -6781 -3282
rect -6777 -3293 -6773 -3282
rect -6828 -3314 -6824 -3294
rect -6820 -3314 -6816 -3294
rect -6650 -3301 -6646 -3290
rect -6642 -3301 -6638 -3290
rect -8098 -3367 -8094 -3347
rect -8090 -3367 -8086 -3347
rect -8066 -3367 -8062 -3347
rect -8058 -3367 -8054 -3347
rect -7829 -3362 -7825 -3342
rect -7821 -3362 -7817 -3342
rect -6693 -3322 -6689 -3302
rect -6685 -3322 -6681 -3302
rect -6502 -3308 -6498 -3298
rect -6494 -3308 -6490 -3298
rect -6566 -3318 -6562 -3308
rect -6558 -3318 -6554 -3308
rect -6533 -3318 -6529 -3308
rect -6525 -3318 -6521 -3308
rect -8195 -3391 -8191 -3371
rect -8187 -3391 -8183 -3371
rect -8143 -3391 -8139 -3371
rect -8135 -3391 -8131 -3371
rect -6340 -3364 -6336 -3354
rect -6332 -3364 -6328 -3354
rect -6404 -3374 -6400 -3364
rect -6396 -3374 -6392 -3364
rect -6371 -3374 -6367 -3364
rect -6363 -3374 -6359 -3364
rect -7786 -3396 -7782 -3385
rect -7778 -3396 -7774 -3385
rect -7829 -3417 -7825 -3397
rect -7821 -3417 -7817 -3397
rect -8299 -3438 -8295 -3418
rect -8291 -3438 -8287 -3418
rect -8247 -3438 -8243 -3418
rect -8239 -3438 -8235 -3418
rect -8195 -3438 -8191 -3418
rect -8187 -3438 -8183 -3418
rect -8143 -3438 -8139 -3418
rect -8135 -3438 -8131 -3418
rect -6182 -3420 -6178 -3410
rect -6174 -3420 -6170 -3410
rect -6246 -3430 -6242 -3420
rect -6238 -3430 -6234 -3420
rect -6213 -3430 -6209 -3420
rect -6205 -3430 -6201 -3420
rect -6016 -3496 -6012 -3486
rect -6008 -3496 -6004 -3486
rect -6080 -3506 -6076 -3496
rect -6072 -3506 -6068 -3496
rect -6047 -3506 -6043 -3496
rect -6039 -3506 -6035 -3496
rect -5712 -3517 -5708 -3497
rect -5704 -3517 -5700 -3497
rect -5680 -3517 -5676 -3497
rect -5672 -3517 -5668 -3497
rect -5809 -3541 -5805 -3521
rect -5801 -3541 -5797 -3521
rect -5757 -3541 -5753 -3521
rect -5749 -3541 -5745 -3521
rect -5545 -3556 -5541 -3545
rect -5537 -3556 -5533 -3545
rect -5913 -3588 -5909 -3568
rect -5905 -3588 -5901 -3568
rect -5861 -3588 -5857 -3568
rect -5853 -3588 -5849 -3568
rect -5809 -3588 -5805 -3568
rect -5801 -3588 -5797 -3568
rect -5757 -3588 -5753 -3568
rect -5749 -3588 -5745 -3568
rect -7864 -3924 -7854 -3920
rect -7864 -3932 -7854 -3928
rect -7764 -3939 -7760 -3931
rect -7756 -3939 -7752 -3931
rect -8043 -3975 -8039 -3955
rect -8035 -3975 -8031 -3955
rect -8011 -3975 -8007 -3955
rect -8003 -3975 -7999 -3955
rect -7864 -3975 -7854 -3971
rect -7764 -3972 -7760 -3962
rect -7756 -3972 -7752 -3962
rect -7728 -3964 -7724 -3954
rect -7720 -3964 -7716 -3954
rect -8140 -3999 -8136 -3979
rect -8132 -3999 -8128 -3979
rect -8088 -3999 -8084 -3979
rect -8080 -3999 -8076 -3979
rect -7864 -3983 -7854 -3979
rect -7603 -4016 -7599 -3996
rect -7595 -4016 -7591 -3996
rect -8244 -4046 -8240 -4026
rect -8236 -4046 -8232 -4026
rect -8192 -4046 -8188 -4026
rect -8184 -4046 -8180 -4026
rect -8140 -4046 -8136 -4026
rect -8132 -4046 -8128 -4026
rect -8088 -4046 -8084 -4026
rect -8080 -4046 -8076 -4026
rect -7434 -4015 -7430 -3995
rect -7426 -4015 -7422 -3995
rect -7270 -4013 -7266 -3993
rect -7262 -4013 -7258 -3993
rect -7130 -4015 -7126 -3995
rect -7122 -4015 -7118 -3995
rect -7560 -4050 -7556 -4039
rect -7552 -4050 -7548 -4039
rect -7391 -4049 -7387 -4038
rect -7383 -4049 -7379 -4038
rect -7227 -4047 -7223 -4036
rect -7219 -4047 -7215 -4036
rect -6979 -4028 -6975 -4008
rect -6971 -4028 -6967 -4008
rect -7603 -4071 -7599 -4051
rect -7595 -4071 -7591 -4051
rect -7434 -4070 -7430 -4050
rect -7426 -4070 -7422 -4050
rect -7270 -4068 -7266 -4048
rect -7262 -4068 -7258 -4048
rect -7087 -4049 -7083 -4038
rect -7079 -4049 -7075 -4038
rect -7130 -4070 -7126 -4050
rect -7122 -4070 -7118 -4050
rect -6936 -4062 -6932 -4051
rect -6928 -4062 -6924 -4051
rect -6639 -4055 -6635 -4045
rect -6631 -4055 -6627 -4045
rect -6979 -4083 -6975 -4063
rect -6971 -4083 -6967 -4063
rect -6703 -4065 -6699 -4055
rect -6695 -4065 -6691 -4055
rect -6670 -4065 -6666 -4055
rect -6662 -4065 -6658 -4055
rect -8026 -4216 -8022 -4196
rect -8018 -4216 -8014 -4196
rect -7994 -4216 -7990 -4196
rect -7986 -4216 -7982 -4196
rect -8123 -4240 -8119 -4220
rect -8115 -4240 -8111 -4220
rect -8071 -4240 -8067 -4220
rect -8063 -4240 -8059 -4220
rect -6816 -4232 -6812 -4212
rect -6808 -4232 -6804 -4212
rect -8227 -4287 -8223 -4267
rect -8219 -4287 -8215 -4267
rect -8175 -4287 -8171 -4267
rect -8167 -4287 -8163 -4267
rect -8123 -4287 -8119 -4267
rect -8115 -4287 -8111 -4267
rect -8071 -4287 -8067 -4267
rect -8063 -4287 -8059 -4267
rect -7836 -4277 -7832 -4257
rect -7828 -4277 -7824 -4257
rect -6773 -4266 -6769 -4255
rect -6765 -4266 -6761 -4255
rect -6505 -4265 -6501 -4255
rect -6497 -4265 -6493 -4255
rect -6816 -4287 -6812 -4267
rect -6808 -4287 -6804 -4267
rect -6569 -4275 -6565 -4265
rect -6561 -4275 -6557 -4265
rect -6536 -4275 -6532 -4265
rect -6528 -4275 -6524 -4265
rect -7793 -4311 -7789 -4300
rect -7785 -4311 -7781 -4300
rect -7836 -4332 -7832 -4312
rect -7828 -4332 -7824 -4312
rect -6197 -4389 -6193 -4385
rect -6189 -4383 -6185 -4379
rect -6358 -4425 -6354 -4415
rect -6350 -4425 -6346 -4415
rect -6422 -4435 -6418 -4425
rect -6414 -4435 -6410 -4425
rect -6389 -4435 -6385 -4425
rect -6381 -4435 -6377 -4425
rect -6197 -4443 -6193 -4439
rect -6189 -4437 -6185 -4433
rect -6179 -4437 -6175 -4433
rect -6171 -4437 -6167 -4433
rect -5879 -4442 -5875 -4422
rect -5871 -4442 -5867 -4422
rect -5847 -4442 -5843 -4422
rect -5839 -4442 -5835 -4422
rect -5976 -4466 -5972 -4446
rect -5968 -4466 -5964 -4446
rect -5924 -4466 -5920 -4446
rect -5916 -4466 -5912 -4446
rect -5721 -4468 -5717 -4457
rect -5713 -4468 -5709 -4457
rect -6080 -4513 -6076 -4493
rect -6072 -4513 -6068 -4493
rect -6028 -4513 -6024 -4493
rect -6020 -4513 -6016 -4493
rect -5976 -4513 -5972 -4493
rect -5968 -4513 -5964 -4493
rect -5924 -4513 -5920 -4493
rect -5916 -4513 -5912 -4493
rect -7864 -4692 -7854 -4688
rect -7864 -4700 -7854 -4696
rect -7764 -4707 -7760 -4699
rect -7756 -4707 -7752 -4699
rect -7864 -4743 -7854 -4739
rect -7764 -4740 -7760 -4730
rect -7756 -4740 -7752 -4730
rect -7728 -4732 -7724 -4722
rect -7720 -4732 -7716 -4722
rect -7864 -4751 -7854 -4747
rect -8037 -4779 -8033 -4759
rect -8029 -4779 -8025 -4759
rect -8005 -4779 -8001 -4759
rect -7997 -4779 -7993 -4759
rect -8134 -4803 -8130 -4783
rect -8126 -4803 -8122 -4783
rect -8082 -4803 -8078 -4783
rect -8074 -4803 -8070 -4783
rect -7582 -4789 -7578 -4769
rect -7574 -4789 -7570 -4769
rect -7539 -4823 -7535 -4812
rect -7531 -4823 -7527 -4812
rect -8238 -4850 -8234 -4830
rect -8230 -4850 -8226 -4830
rect -8186 -4850 -8182 -4830
rect -8178 -4850 -8174 -4830
rect -8134 -4850 -8130 -4830
rect -8126 -4850 -8122 -4830
rect -8082 -4850 -8078 -4830
rect -8074 -4850 -8070 -4830
rect -7582 -4844 -7578 -4824
rect -7574 -4844 -7570 -4824
rect -7386 -4915 -7382 -4905
rect -7378 -4915 -7374 -4905
rect -7450 -4925 -7446 -4915
rect -7442 -4925 -7438 -4915
rect -7417 -4925 -7413 -4915
rect -7409 -4925 -7405 -4915
rect -7581 -4994 -7577 -4974
rect -7573 -4994 -7569 -4974
rect -7538 -5028 -7534 -5017
rect -7530 -5028 -7526 -5017
rect -7115 -5000 -7111 -4996
rect -7107 -4994 -7103 -4990
rect -7240 -5028 -7236 -5018
rect -7232 -5028 -7228 -5018
rect -7581 -5049 -7577 -5029
rect -7573 -5049 -7569 -5029
rect -7304 -5038 -7300 -5028
rect -7296 -5038 -7292 -5028
rect -7271 -5038 -7267 -5028
rect -7263 -5038 -7259 -5028
rect -8024 -5091 -8020 -5071
rect -8016 -5091 -8012 -5071
rect -7992 -5091 -7988 -5071
rect -7984 -5091 -7980 -5071
rect -7115 -5054 -7111 -5050
rect -7107 -5048 -7103 -5044
rect -7097 -5048 -7093 -5044
rect -7089 -5048 -7085 -5044
rect -8121 -5115 -8117 -5095
rect -8113 -5115 -8109 -5095
rect -8069 -5115 -8065 -5095
rect -8061 -5115 -8057 -5095
rect -6798 -5051 -6794 -5031
rect -6790 -5051 -6786 -5031
rect -6766 -5051 -6762 -5031
rect -6758 -5051 -6754 -5031
rect -6895 -5075 -6891 -5055
rect -6887 -5075 -6883 -5055
rect -6843 -5075 -6839 -5055
rect -6835 -5075 -6831 -5055
rect -7842 -5126 -7838 -5106
rect -7834 -5126 -7830 -5106
rect -6687 -5088 -6683 -5077
rect -6679 -5088 -6675 -5077
rect -3990 -5100 -3986 -5096
rect -3982 -5094 -3978 -5090
rect -6999 -5122 -6995 -5102
rect -6991 -5122 -6987 -5102
rect -6947 -5122 -6943 -5102
rect -6939 -5122 -6935 -5102
rect -6895 -5122 -6891 -5102
rect -6887 -5122 -6883 -5102
rect -6843 -5122 -6839 -5102
rect -6835 -5122 -6831 -5102
rect -8225 -5162 -8221 -5142
rect -8217 -5162 -8213 -5142
rect -8173 -5162 -8169 -5142
rect -8165 -5162 -8161 -5142
rect -8121 -5162 -8117 -5142
rect -8113 -5162 -8109 -5142
rect -8069 -5162 -8065 -5142
rect -8061 -5162 -8057 -5142
rect -7799 -5160 -7795 -5149
rect -7791 -5160 -7787 -5149
rect -3990 -5154 -3986 -5150
rect -3982 -5148 -3978 -5144
rect -3972 -5148 -3968 -5144
rect -3964 -5148 -3960 -5144
rect -7842 -5181 -7838 -5161
rect -7834 -5181 -7830 -5161
rect -7886 -5454 -7876 -5450
rect -7886 -5462 -7876 -5458
rect -8037 -5485 -8033 -5465
rect -8029 -5485 -8025 -5465
rect -8005 -5485 -8001 -5465
rect -7997 -5485 -7993 -5465
rect -7786 -5469 -7782 -5461
rect -7778 -5469 -7774 -5461
rect -8134 -5509 -8130 -5489
rect -8126 -5509 -8122 -5489
rect -8082 -5509 -8078 -5489
rect -8074 -5509 -8070 -5489
rect -7886 -5505 -7876 -5501
rect -7786 -5502 -7782 -5492
rect -7778 -5502 -7774 -5492
rect -7750 -5494 -7746 -5484
rect -7742 -5494 -7738 -5484
rect -7886 -5513 -7876 -5509
rect -8238 -5556 -8234 -5536
rect -8230 -5556 -8226 -5536
rect -8186 -5556 -8182 -5536
rect -8178 -5556 -8174 -5536
rect -8134 -5556 -8130 -5536
rect -8126 -5556 -8122 -5536
rect -8082 -5556 -8078 -5536
rect -8074 -5556 -8070 -5536
rect -7670 -5569 -7666 -5549
rect -7662 -5569 -7658 -5549
rect -7627 -5603 -7623 -5592
rect -7619 -5603 -7615 -5592
rect -7670 -5624 -7666 -5604
rect -7662 -5624 -7658 -5604
rect -8034 -5734 -8030 -5714
rect -8026 -5734 -8022 -5714
rect -8002 -5734 -7998 -5714
rect -7994 -5734 -7990 -5714
rect -8131 -5758 -8127 -5738
rect -8123 -5758 -8119 -5738
rect -8079 -5758 -8075 -5738
rect -8071 -5758 -8067 -5738
rect -7839 -5749 -7835 -5729
rect -7831 -5749 -7827 -5729
rect -7307 -5724 -7303 -5720
rect -7299 -5718 -7295 -5714
rect -6982 -5705 -6978 -5685
rect -6974 -5705 -6970 -5685
rect -6950 -5705 -6946 -5685
rect -6942 -5705 -6938 -5685
rect -7079 -5729 -7075 -5709
rect -7071 -5729 -7067 -5709
rect -7027 -5729 -7023 -5709
rect -7019 -5729 -7015 -5709
rect -7492 -5758 -7488 -5748
rect -7484 -5758 -7480 -5748
rect -7556 -5768 -7552 -5758
rect -7548 -5768 -7544 -5758
rect -7523 -5768 -7519 -5758
rect -7515 -5768 -7511 -5758
rect -7796 -5783 -7792 -5772
rect -7788 -5783 -7784 -5772
rect -7307 -5778 -7303 -5774
rect -7299 -5772 -7295 -5768
rect -7289 -5772 -7285 -5768
rect -7281 -5772 -7277 -5768
rect -7183 -5776 -7179 -5756
rect -7175 -5776 -7171 -5756
rect -7131 -5776 -7127 -5756
rect -7123 -5776 -7119 -5756
rect -7079 -5776 -7075 -5756
rect -7071 -5776 -7067 -5756
rect -7027 -5776 -7023 -5756
rect -7019 -5776 -7015 -5756
rect -6823 -5763 -6819 -5752
rect -6815 -5763 -6811 -5752
rect -8235 -5805 -8231 -5785
rect -8227 -5805 -8223 -5785
rect -8183 -5805 -8179 -5785
rect -8175 -5805 -8171 -5785
rect -8131 -5805 -8127 -5785
rect -8123 -5805 -8119 -5785
rect -8079 -5805 -8075 -5785
rect -8071 -5805 -8067 -5785
rect -7839 -5804 -7835 -5784
rect -7831 -5804 -7827 -5784
rect -7635 -5840 -7631 -5836
rect -7627 -5834 -7623 -5830
rect -7635 -5894 -7631 -5890
rect -7627 -5888 -7623 -5884
rect -7617 -5888 -7613 -5884
rect -7609 -5888 -7605 -5884
rect -7259 -5945 -7255 -5925
rect -7251 -5945 -7247 -5925
rect -7227 -5945 -7223 -5925
rect -7219 -5945 -7215 -5925
rect -7356 -5969 -7352 -5949
rect -7348 -5969 -7344 -5949
rect -7304 -5969 -7300 -5949
rect -7296 -5969 -7292 -5949
rect -7124 -5985 -7120 -5974
rect -7116 -5985 -7112 -5974
rect -7460 -6016 -7456 -5996
rect -7452 -6016 -7448 -5996
rect -7408 -6016 -7404 -5996
rect -7400 -6016 -7396 -5996
rect -7356 -6016 -7352 -5996
rect -7348 -6016 -7344 -5996
rect -7304 -6016 -7300 -5996
rect -7296 -6016 -7292 -5996
rect -7659 -6045 -7655 -6025
rect -7651 -6045 -7647 -6025
rect -7627 -6045 -7623 -6025
rect -7619 -6045 -7615 -6025
rect -7756 -6069 -7752 -6049
rect -7748 -6069 -7744 -6049
rect -7704 -6069 -7700 -6049
rect -7696 -6069 -7692 -6049
rect -7860 -6116 -7856 -6096
rect -7852 -6116 -7848 -6096
rect -7808 -6116 -7804 -6096
rect -7800 -6116 -7796 -6096
rect -7756 -6116 -7752 -6096
rect -7748 -6116 -7744 -6096
rect -7704 -6116 -7700 -6096
rect -7696 -6116 -7692 -6096
rect -7548 -6230 -7544 -6219
rect -7540 -6230 -7536 -6219
<< pdcontact >>
rect -2918 -530 -2914 -510
rect -2910 -530 -2906 -510
rect -2891 -530 -2887 -510
rect -2883 -530 -2879 -510
rect -2856 -600 -2852 -560
rect -2848 -600 -2844 -560
rect -2540 -600 -2520 -596
rect -2540 -608 -2520 -604
rect -2442 -612 -2438 -592
rect -2434 -612 -2430 -592
rect -2540 -651 -2520 -647
rect -2540 -659 -2520 -655
rect -2288 -678 -2284 -658
rect -2280 -678 -2276 -658
rect -2288 -725 -2284 -706
rect -2280 -725 -2276 -706
rect -2239 -722 -2235 -702
rect -2231 -722 -2227 -702
rect -1990 -708 -1986 -668
rect -1982 -708 -1978 -668
rect -1938 -708 -1934 -668
rect -1930 -708 -1926 -668
rect -1886 -708 -1882 -668
rect -1878 -708 -1874 -668
rect -1834 -708 -1830 -668
rect -1826 -708 -1822 -668
rect -1789 -700 -1785 -660
rect -1781 -700 -1777 -660
rect -1757 -700 -1753 -660
rect -1749 -700 -1745 -660
rect -1990 -770 -1986 -730
rect -1982 -770 -1978 -730
rect -1938 -770 -1934 -730
rect -1930 -770 -1926 -730
rect -8313 -3031 -8309 -2991
rect -8305 -3031 -8301 -2991
rect -8261 -3031 -8257 -2991
rect -8253 -3031 -8249 -2991
rect -8209 -3031 -8205 -2991
rect -8201 -3031 -8197 -2991
rect -8157 -3031 -8153 -2991
rect -8149 -3031 -8145 -2991
rect -8112 -3023 -8108 -2983
rect -8104 -3023 -8100 -2983
rect -8080 -3023 -8076 -2983
rect -8072 -3023 -8068 -2983
rect -8313 -3093 -8309 -3053
rect -8305 -3093 -8301 -3053
rect -8261 -3093 -8257 -3053
rect -8253 -3093 -8249 -3053
rect -7832 -3073 -7812 -3069
rect -7832 -3081 -7812 -3077
rect -7734 -3085 -7730 -3065
rect -7726 -3085 -7722 -3065
rect -7832 -3124 -7812 -3120
rect -7630 -3127 -7626 -3107
rect -7622 -3127 -7618 -3107
rect -7603 -3127 -7599 -3107
rect -7595 -3127 -7591 -3107
rect -7832 -3132 -7812 -3128
rect -7568 -3197 -7564 -3157
rect -7560 -3197 -7556 -3157
rect -7485 -3165 -7481 -3145
rect -7477 -3165 -7473 -3145
rect -7458 -3165 -7454 -3145
rect -7450 -3165 -7446 -3145
rect -7292 -3181 -7288 -3161
rect -7284 -3181 -7280 -3161
rect -7265 -3181 -7261 -3161
rect -7257 -3181 -7253 -3161
rect -7146 -3179 -7142 -3159
rect -7138 -3179 -7134 -3159
rect -7119 -3179 -7115 -3159
rect -7111 -3179 -7107 -3159
rect -7423 -3235 -7419 -3195
rect -7415 -3235 -7411 -3195
rect -7002 -3183 -6998 -3163
rect -6994 -3183 -6990 -3163
rect -6975 -3183 -6971 -3163
rect -6967 -3183 -6963 -3163
rect -7230 -3251 -7226 -3211
rect -7222 -3251 -7218 -3211
rect -6847 -3185 -6843 -3165
rect -6839 -3185 -6835 -3165
rect -6820 -3185 -6816 -3165
rect -6812 -3185 -6808 -3165
rect -8299 -3335 -8295 -3295
rect -8291 -3335 -8287 -3295
rect -8247 -3335 -8243 -3295
rect -8239 -3335 -8235 -3295
rect -8195 -3335 -8191 -3295
rect -8187 -3335 -8183 -3295
rect -8143 -3335 -8139 -3295
rect -8135 -3335 -8131 -3295
rect -8098 -3327 -8094 -3287
rect -8090 -3327 -8086 -3287
rect -8066 -3327 -8062 -3287
rect -8058 -3327 -8054 -3287
rect -7848 -3288 -7844 -3268
rect -7840 -3288 -7836 -3268
rect -7821 -3288 -7817 -3268
rect -7813 -3288 -7809 -3268
rect -7084 -3249 -7080 -3209
rect -7076 -3249 -7072 -3209
rect -6712 -3193 -6708 -3173
rect -6704 -3193 -6700 -3173
rect -6685 -3193 -6681 -3173
rect -6677 -3193 -6673 -3173
rect -6940 -3253 -6936 -3213
rect -6932 -3253 -6928 -3213
rect -6785 -3255 -6781 -3215
rect -6777 -3255 -6773 -3215
rect -6650 -3263 -6646 -3223
rect -6642 -3263 -6638 -3223
rect -6551 -3236 -6547 -3216
rect -6543 -3236 -6539 -3216
rect -6551 -3283 -6547 -3264
rect -6543 -3283 -6539 -3264
rect -8299 -3397 -8295 -3357
rect -8291 -3397 -8287 -3357
rect -8247 -3397 -8243 -3357
rect -8239 -3397 -8235 -3357
rect -7786 -3358 -7782 -3318
rect -7778 -3358 -7774 -3318
rect -6502 -3280 -6498 -3260
rect -6494 -3280 -6490 -3260
rect -6389 -3292 -6385 -3272
rect -6381 -3292 -6377 -3272
rect -6389 -3339 -6385 -3320
rect -6381 -3339 -6377 -3320
rect -6340 -3336 -6336 -3316
rect -6332 -3336 -6328 -3316
rect -6231 -3348 -6227 -3328
rect -6223 -3348 -6219 -3328
rect -6231 -3395 -6227 -3376
rect -6223 -3395 -6219 -3376
rect -6182 -3392 -6178 -3372
rect -6174 -3392 -6170 -3372
rect -6065 -3424 -6061 -3404
rect -6057 -3424 -6053 -3404
rect -6065 -3471 -6061 -3452
rect -6057 -3471 -6053 -3452
rect -6016 -3468 -6012 -3448
rect -6008 -3468 -6004 -3448
rect -5913 -3485 -5909 -3445
rect -5905 -3485 -5901 -3445
rect -5861 -3485 -5857 -3445
rect -5853 -3485 -5849 -3445
rect -5809 -3485 -5805 -3445
rect -5801 -3485 -5797 -3445
rect -5757 -3485 -5753 -3445
rect -5749 -3485 -5745 -3445
rect -5712 -3477 -5708 -3437
rect -5704 -3477 -5700 -3437
rect -5680 -3477 -5676 -3437
rect -5672 -3477 -5668 -3437
rect -5913 -3547 -5909 -3507
rect -5905 -3547 -5901 -3507
rect -5861 -3547 -5857 -3507
rect -5853 -3547 -5849 -3507
rect -5545 -3518 -5541 -3478
rect -5537 -3518 -5533 -3478
rect -8244 -3943 -8240 -3903
rect -8236 -3943 -8232 -3903
rect -8192 -3943 -8188 -3903
rect -8184 -3943 -8180 -3903
rect -8140 -3943 -8136 -3903
rect -8132 -3943 -8128 -3903
rect -8088 -3943 -8084 -3903
rect -8080 -3943 -8076 -3903
rect -8043 -3935 -8039 -3895
rect -8035 -3935 -8031 -3895
rect -8011 -3935 -8007 -3895
rect -8003 -3935 -7999 -3895
rect -7826 -3924 -7806 -3920
rect -7826 -3932 -7806 -3928
rect -7728 -3936 -7724 -3916
rect -7720 -3936 -7716 -3916
rect -8244 -4005 -8240 -3965
rect -8236 -4005 -8232 -3965
rect -8192 -4005 -8188 -3965
rect -8184 -4005 -8180 -3965
rect -7622 -3942 -7618 -3922
rect -7614 -3942 -7610 -3922
rect -7595 -3942 -7591 -3922
rect -7587 -3942 -7583 -3922
rect -7453 -3941 -7449 -3921
rect -7445 -3941 -7441 -3921
rect -7426 -3941 -7422 -3921
rect -7418 -3941 -7414 -3921
rect -7289 -3939 -7285 -3919
rect -7281 -3939 -7277 -3919
rect -7262 -3939 -7258 -3919
rect -7254 -3939 -7250 -3919
rect -7826 -3975 -7806 -3971
rect -7149 -3941 -7145 -3921
rect -7141 -3941 -7137 -3921
rect -7122 -3941 -7118 -3921
rect -7114 -3941 -7110 -3921
rect -6998 -3954 -6994 -3934
rect -6990 -3954 -6986 -3934
rect -6971 -3954 -6967 -3934
rect -6963 -3954 -6959 -3934
rect -7826 -3983 -7806 -3979
rect -7560 -4012 -7556 -3972
rect -7552 -4012 -7548 -3972
rect -7391 -4011 -7387 -3971
rect -7383 -4011 -7379 -3971
rect -7227 -4009 -7223 -3969
rect -7219 -4009 -7215 -3969
rect -7087 -4011 -7083 -3971
rect -7079 -4011 -7075 -3971
rect -6688 -3983 -6684 -3963
rect -6680 -3983 -6676 -3963
rect -6936 -4024 -6932 -3984
rect -6928 -4024 -6924 -3984
rect -6688 -4030 -6684 -4011
rect -6680 -4030 -6676 -4011
rect -6639 -4027 -6635 -4007
rect -6631 -4027 -6627 -4007
rect -8227 -4184 -8223 -4144
rect -8219 -4184 -8215 -4144
rect -8175 -4184 -8171 -4144
rect -8167 -4184 -8163 -4144
rect -8123 -4184 -8119 -4144
rect -8115 -4184 -8111 -4144
rect -8071 -4184 -8067 -4144
rect -8063 -4184 -8059 -4144
rect -8026 -4176 -8022 -4136
rect -8018 -4176 -8014 -4136
rect -7994 -4176 -7990 -4136
rect -7986 -4176 -7982 -4136
rect -6835 -4158 -6831 -4138
rect -6827 -4158 -6823 -4138
rect -6808 -4158 -6804 -4138
rect -6800 -4158 -6796 -4138
rect -8227 -4246 -8223 -4206
rect -8219 -4246 -8215 -4206
rect -8175 -4246 -8171 -4206
rect -8167 -4246 -8163 -4206
rect -7855 -4203 -7851 -4183
rect -7847 -4203 -7843 -4183
rect -7828 -4203 -7824 -4183
rect -7820 -4203 -7816 -4183
rect -6773 -4228 -6769 -4188
rect -6765 -4228 -6761 -4188
rect -6554 -4193 -6550 -4173
rect -6546 -4193 -6542 -4173
rect -7793 -4273 -7789 -4233
rect -7785 -4273 -7781 -4233
rect -6554 -4240 -6550 -4221
rect -6546 -4240 -6542 -4221
rect -6505 -4237 -6501 -4217
rect -6497 -4237 -6493 -4217
rect -6407 -4353 -6403 -4333
rect -6399 -4353 -6395 -4333
rect -6197 -4350 -6193 -4346
rect -6407 -4400 -6403 -4381
rect -6399 -4400 -6395 -4381
rect -6189 -4366 -6185 -4362
rect -6358 -4397 -6354 -4377
rect -6350 -4397 -6346 -4377
rect -6197 -4405 -6193 -4401
rect -6189 -4421 -6185 -4417
rect -6179 -4421 -6175 -4417
rect -6080 -4410 -6076 -4370
rect -6072 -4410 -6068 -4370
rect -6028 -4410 -6024 -4370
rect -6020 -4410 -6016 -4370
rect -5976 -4410 -5972 -4370
rect -5968 -4410 -5964 -4370
rect -5924 -4410 -5920 -4370
rect -5916 -4410 -5912 -4370
rect -5879 -4402 -5875 -4362
rect -5871 -4402 -5867 -4362
rect -5847 -4402 -5843 -4362
rect -5839 -4402 -5835 -4362
rect -6171 -4421 -6167 -4417
rect -6080 -4472 -6076 -4432
rect -6072 -4472 -6068 -4432
rect -6028 -4472 -6024 -4432
rect -6020 -4472 -6016 -4432
rect -5721 -4430 -5717 -4390
rect -5713 -4430 -5709 -4390
rect -7826 -4692 -7806 -4688
rect -8238 -4747 -8234 -4707
rect -8230 -4747 -8226 -4707
rect -8186 -4747 -8182 -4707
rect -8178 -4747 -8174 -4707
rect -8134 -4747 -8130 -4707
rect -8126 -4747 -8122 -4707
rect -8082 -4747 -8078 -4707
rect -8074 -4747 -8070 -4707
rect -8037 -4739 -8033 -4699
rect -8029 -4739 -8025 -4699
rect -8005 -4739 -8001 -4699
rect -7997 -4739 -7993 -4699
rect -7826 -4700 -7806 -4696
rect -7728 -4704 -7724 -4684
rect -7720 -4704 -7716 -4684
rect -7601 -4715 -7597 -4695
rect -7593 -4715 -7589 -4695
rect -7574 -4715 -7570 -4695
rect -7566 -4715 -7562 -4695
rect -7826 -4743 -7806 -4739
rect -7826 -4751 -7806 -4747
rect -8238 -4809 -8234 -4769
rect -8230 -4809 -8226 -4769
rect -8186 -4809 -8182 -4769
rect -8178 -4809 -8174 -4769
rect -7539 -4785 -7535 -4745
rect -7531 -4785 -7527 -4745
rect -7435 -4843 -7431 -4823
rect -7427 -4843 -7423 -4823
rect -7435 -4890 -7431 -4871
rect -7427 -4890 -7423 -4871
rect -7600 -4920 -7596 -4900
rect -7592 -4920 -7588 -4900
rect -7573 -4920 -7569 -4900
rect -7565 -4920 -7561 -4900
rect -7386 -4887 -7382 -4867
rect -7378 -4887 -7374 -4867
rect -7538 -4990 -7534 -4950
rect -7530 -4990 -7526 -4950
rect -7289 -4956 -7285 -4936
rect -7281 -4956 -7277 -4936
rect -7115 -4961 -7111 -4957
rect -8225 -5059 -8221 -5019
rect -8217 -5059 -8213 -5019
rect -8173 -5059 -8169 -5019
rect -8165 -5059 -8161 -5019
rect -8121 -5059 -8117 -5019
rect -8113 -5059 -8109 -5019
rect -8069 -5059 -8065 -5019
rect -8061 -5059 -8057 -5019
rect -8024 -5051 -8020 -5011
rect -8016 -5051 -8012 -5011
rect -7992 -5051 -7988 -5011
rect -7984 -5051 -7980 -5011
rect -7289 -5003 -7285 -4984
rect -7281 -5003 -7277 -4984
rect -7107 -4977 -7103 -4973
rect -7240 -5000 -7236 -4980
rect -7232 -5000 -7228 -4980
rect -7115 -5016 -7111 -5012
rect -7861 -5052 -7857 -5032
rect -7853 -5052 -7849 -5032
rect -7834 -5052 -7830 -5032
rect -7826 -5052 -7822 -5032
rect -7107 -5032 -7103 -5028
rect -7097 -5032 -7093 -5028
rect -6999 -5019 -6995 -4979
rect -6991 -5019 -6987 -4979
rect -6947 -5019 -6943 -4979
rect -6939 -5019 -6935 -4979
rect -6895 -5019 -6891 -4979
rect -6887 -5019 -6883 -4979
rect -6843 -5019 -6839 -4979
rect -6835 -5019 -6831 -4979
rect -6798 -5011 -6794 -4971
rect -6790 -5011 -6786 -4971
rect -6766 -5011 -6762 -4971
rect -6758 -5011 -6754 -4971
rect -7089 -5032 -7085 -5028
rect -8225 -5121 -8221 -5081
rect -8217 -5121 -8213 -5081
rect -8173 -5121 -8169 -5081
rect -8165 -5121 -8161 -5081
rect -6999 -5081 -6995 -5041
rect -6991 -5081 -6987 -5041
rect -6947 -5081 -6943 -5041
rect -6939 -5081 -6935 -5041
rect -6687 -5050 -6683 -5010
rect -6679 -5050 -6675 -5010
rect -3990 -5061 -3986 -5057
rect -3982 -5077 -3978 -5073
rect -7799 -5122 -7795 -5082
rect -7791 -5122 -7787 -5082
rect -3990 -5116 -3986 -5112
rect -3982 -5132 -3978 -5128
rect -3972 -5132 -3968 -5128
rect -3964 -5132 -3960 -5128
rect -8238 -5453 -8234 -5413
rect -8230 -5453 -8226 -5413
rect -8186 -5453 -8182 -5413
rect -8178 -5453 -8174 -5413
rect -8134 -5453 -8130 -5413
rect -8126 -5453 -8122 -5413
rect -8082 -5453 -8078 -5413
rect -8074 -5453 -8070 -5413
rect -8037 -5445 -8033 -5405
rect -8029 -5445 -8025 -5405
rect -8005 -5445 -8001 -5405
rect -7997 -5445 -7993 -5405
rect -7848 -5454 -7828 -5450
rect -7848 -5462 -7828 -5458
rect -8238 -5515 -8234 -5475
rect -8230 -5515 -8226 -5475
rect -8186 -5515 -8182 -5475
rect -8178 -5515 -8174 -5475
rect -7750 -5466 -7746 -5446
rect -7742 -5466 -7738 -5446
rect -7848 -5505 -7828 -5501
rect -7689 -5495 -7685 -5475
rect -7681 -5495 -7677 -5475
rect -7662 -5495 -7658 -5475
rect -7654 -5495 -7650 -5475
rect -7848 -5513 -7828 -5509
rect -7627 -5565 -7623 -5525
rect -7619 -5565 -7615 -5525
rect -8235 -5702 -8231 -5662
rect -8227 -5702 -8223 -5662
rect -8183 -5702 -8179 -5662
rect -8175 -5702 -8171 -5662
rect -8131 -5702 -8127 -5662
rect -8123 -5702 -8119 -5662
rect -8079 -5702 -8075 -5662
rect -8071 -5702 -8067 -5662
rect -8034 -5694 -8030 -5654
rect -8026 -5694 -8022 -5654
rect -8002 -5694 -7998 -5654
rect -7994 -5694 -7990 -5654
rect -7858 -5675 -7854 -5655
rect -7850 -5675 -7846 -5655
rect -7831 -5675 -7827 -5655
rect -7823 -5675 -7819 -5655
rect -7541 -5686 -7537 -5666
rect -7533 -5686 -7529 -5666
rect -7183 -5673 -7179 -5633
rect -7175 -5673 -7171 -5633
rect -7131 -5673 -7127 -5633
rect -7123 -5673 -7119 -5633
rect -7079 -5673 -7075 -5633
rect -7071 -5673 -7067 -5633
rect -7027 -5673 -7023 -5633
rect -7019 -5673 -7015 -5633
rect -6982 -5665 -6978 -5625
rect -6974 -5665 -6970 -5625
rect -6950 -5665 -6946 -5625
rect -6942 -5665 -6938 -5625
rect -7307 -5685 -7303 -5681
rect -8235 -5764 -8231 -5724
rect -8227 -5764 -8223 -5724
rect -8183 -5764 -8179 -5724
rect -8175 -5764 -8171 -5724
rect -7796 -5745 -7792 -5705
rect -7788 -5745 -7784 -5705
rect -7541 -5733 -7537 -5714
rect -7533 -5733 -7529 -5714
rect -7299 -5701 -7295 -5697
rect -7492 -5730 -7488 -5710
rect -7484 -5730 -7480 -5710
rect -7183 -5735 -7179 -5695
rect -7175 -5735 -7171 -5695
rect -7131 -5735 -7127 -5695
rect -7123 -5735 -7119 -5695
rect -6823 -5725 -6819 -5685
rect -6815 -5725 -6811 -5685
rect -7307 -5740 -7303 -5736
rect -7299 -5756 -7295 -5752
rect -7289 -5756 -7285 -5752
rect -7281 -5756 -7277 -5752
rect -7635 -5801 -7631 -5797
rect -7627 -5817 -7623 -5813
rect -7635 -5856 -7631 -5852
rect -7627 -5872 -7623 -5868
rect -7617 -5872 -7613 -5868
rect -7609 -5872 -7605 -5868
rect -7460 -5913 -7456 -5873
rect -7452 -5913 -7448 -5873
rect -7408 -5913 -7404 -5873
rect -7400 -5913 -7396 -5873
rect -7356 -5913 -7352 -5873
rect -7348 -5913 -7344 -5873
rect -7304 -5913 -7300 -5873
rect -7296 -5913 -7292 -5873
rect -7259 -5905 -7255 -5865
rect -7251 -5905 -7247 -5865
rect -7227 -5905 -7223 -5865
rect -7219 -5905 -7215 -5865
rect -7860 -6013 -7856 -5973
rect -7852 -6013 -7848 -5973
rect -7808 -6013 -7804 -5973
rect -7800 -6013 -7796 -5973
rect -7756 -6013 -7752 -5973
rect -7748 -6013 -7744 -5973
rect -7704 -6013 -7700 -5973
rect -7696 -6013 -7692 -5973
rect -7659 -6005 -7655 -5965
rect -7651 -6005 -7647 -5965
rect -7627 -6005 -7623 -5965
rect -7619 -6005 -7615 -5965
rect -7460 -5975 -7456 -5935
rect -7452 -5975 -7448 -5935
rect -7408 -5975 -7404 -5935
rect -7400 -5975 -7396 -5935
rect -7124 -5947 -7120 -5907
rect -7116 -5947 -7112 -5907
rect -7860 -6075 -7856 -6035
rect -7852 -6075 -7848 -6035
rect -7808 -6075 -7804 -6035
rect -7800 -6075 -7796 -6035
rect -7548 -6192 -7544 -6152
rect -7540 -6192 -7536 -6152
<< psubstratepcontact >>
rect -2589 -593 -2585 -589
rect -2589 -614 -2585 -610
rect -2589 -644 -2585 -640
rect -2863 -649 -2859 -645
rect -2842 -649 -2838 -645
rect -2449 -655 -2445 -651
rect -2428 -655 -2424 -651
rect -2589 -665 -2585 -661
rect -2906 -670 -2902 -666
rect -2885 -670 -2881 -666
rect -2246 -765 -2242 -761
rect -2225 -765 -2221 -761
rect -2310 -772 -2306 -768
rect -2289 -772 -2285 -768
rect -2277 -772 -2273 -768
rect -2256 -772 -2252 -768
rect -1797 -753 -1793 -749
rect -1773 -753 -1769 -749
rect -1765 -753 -1761 -749
rect -1741 -753 -1737 -749
rect -1973 -824 -1969 -820
rect -1921 -824 -1917 -820
rect -1869 -824 -1865 -820
rect -1817 -824 -1813 -820
rect -7881 -3066 -7877 -3062
rect -8120 -3076 -8116 -3072
rect -8096 -3076 -8092 -3072
rect -8088 -3076 -8084 -3072
rect -8064 -3076 -8060 -3072
rect -7881 -3087 -7877 -3083
rect -7881 -3117 -7877 -3113
rect -7741 -3128 -7737 -3124
rect -7720 -3128 -7716 -3124
rect -7881 -3138 -7877 -3134
rect -8296 -3147 -8292 -3143
rect -8244 -3147 -8240 -3143
rect -8192 -3147 -8188 -3143
rect -8140 -3147 -8136 -3143
rect -7575 -3246 -7571 -3242
rect -7554 -3246 -7550 -3242
rect -7618 -3267 -7614 -3263
rect -7597 -3267 -7593 -3263
rect -7430 -3284 -7426 -3280
rect -7409 -3284 -7405 -3280
rect -7473 -3305 -7469 -3301
rect -7452 -3305 -7448 -3301
rect -7237 -3300 -7233 -3296
rect -7216 -3300 -7212 -3296
rect -7091 -3298 -7087 -3294
rect -7070 -3298 -7066 -3294
rect -6947 -3302 -6943 -3298
rect -6926 -3302 -6922 -3298
rect -6792 -3304 -6788 -3300
rect -6771 -3304 -6767 -3300
rect -7280 -3321 -7276 -3317
rect -7259 -3321 -7255 -3317
rect -7134 -3319 -7130 -3315
rect -7113 -3319 -7109 -3315
rect -6990 -3323 -6986 -3319
rect -6969 -3323 -6965 -3319
rect -6835 -3325 -6831 -3321
rect -6814 -3325 -6810 -3321
rect -6657 -3312 -6653 -3308
rect -6636 -3312 -6632 -3308
rect -6509 -3323 -6505 -3319
rect -6488 -3323 -6484 -3319
rect -6700 -3333 -6696 -3329
rect -6679 -3333 -6675 -3329
rect -6573 -3330 -6569 -3326
rect -6552 -3330 -6548 -3326
rect -6540 -3330 -6536 -3326
rect -6519 -3330 -6515 -3326
rect -8106 -3380 -8102 -3376
rect -8082 -3380 -8078 -3376
rect -8074 -3380 -8070 -3376
rect -8050 -3380 -8046 -3376
rect -6347 -3379 -6343 -3375
rect -6326 -3379 -6322 -3375
rect -6411 -3386 -6407 -3382
rect -6390 -3386 -6386 -3382
rect -6378 -3386 -6374 -3382
rect -6357 -3386 -6353 -3382
rect -7793 -3407 -7789 -3403
rect -7772 -3407 -7768 -3403
rect -7836 -3428 -7832 -3424
rect -7815 -3428 -7811 -3424
rect -6189 -3435 -6185 -3431
rect -6168 -3435 -6164 -3431
rect -6253 -3442 -6249 -3438
rect -6232 -3442 -6228 -3438
rect -6220 -3442 -6216 -3438
rect -6199 -3442 -6195 -3438
rect -8282 -3451 -8278 -3447
rect -8230 -3451 -8226 -3447
rect -8178 -3451 -8174 -3447
rect -8126 -3451 -8122 -3447
rect -6023 -3511 -6019 -3507
rect -6002 -3511 -5998 -3507
rect -6087 -3518 -6083 -3514
rect -6066 -3518 -6062 -3514
rect -6054 -3518 -6050 -3514
rect -6033 -3518 -6029 -3514
rect -5720 -3530 -5716 -3526
rect -5696 -3530 -5692 -3526
rect -5688 -3530 -5684 -3526
rect -5664 -3530 -5660 -3526
rect -5552 -3567 -5548 -3563
rect -5531 -3567 -5527 -3563
rect -5896 -3601 -5892 -3597
rect -5844 -3601 -5840 -3597
rect -5792 -3601 -5788 -3597
rect -5740 -3601 -5736 -3597
rect -7875 -3917 -7871 -3913
rect -7875 -3938 -7871 -3934
rect -7875 -3968 -7871 -3964
rect -7735 -3979 -7731 -3975
rect -7714 -3979 -7710 -3975
rect -8051 -3988 -8047 -3984
rect -8027 -3988 -8023 -3984
rect -8019 -3988 -8015 -3984
rect -7995 -3988 -7991 -3984
rect -7875 -3989 -7871 -3985
rect -8227 -4059 -8223 -4055
rect -8175 -4059 -8171 -4055
rect -8123 -4059 -8119 -4055
rect -8071 -4059 -8067 -4055
rect -7567 -4061 -7563 -4057
rect -7546 -4061 -7542 -4057
rect -7398 -4060 -7394 -4056
rect -7377 -4060 -7373 -4056
rect -7234 -4058 -7230 -4054
rect -7213 -4058 -7209 -4054
rect -7094 -4060 -7090 -4056
rect -7073 -4060 -7069 -4056
rect -7610 -4082 -7606 -4078
rect -7589 -4082 -7585 -4078
rect -7441 -4081 -7437 -4077
rect -7420 -4081 -7416 -4077
rect -7277 -4079 -7273 -4075
rect -7256 -4079 -7252 -4075
rect -7137 -4081 -7133 -4077
rect -7116 -4081 -7112 -4077
rect -6943 -4073 -6939 -4069
rect -6922 -4073 -6918 -4069
rect -6646 -4070 -6642 -4066
rect -6625 -4070 -6621 -4066
rect -6710 -4077 -6706 -4073
rect -6689 -4077 -6685 -4073
rect -6677 -4077 -6673 -4073
rect -6656 -4077 -6652 -4073
rect -6986 -4094 -6982 -4090
rect -6965 -4094 -6961 -4090
rect -8034 -4229 -8030 -4225
rect -8010 -4229 -8006 -4225
rect -8002 -4229 -7998 -4225
rect -7978 -4229 -7974 -4225
rect -8210 -4300 -8206 -4296
rect -8158 -4300 -8154 -4296
rect -8106 -4300 -8102 -4296
rect -8054 -4300 -8050 -4296
rect -6780 -4277 -6776 -4273
rect -6759 -4277 -6755 -4273
rect -6512 -4280 -6508 -4276
rect -6491 -4280 -6487 -4276
rect -6576 -4287 -6572 -4283
rect -6555 -4287 -6551 -4283
rect -6543 -4287 -6539 -4283
rect -6522 -4287 -6518 -4283
rect -6823 -4298 -6819 -4294
rect -6802 -4298 -6798 -4294
rect -7800 -4322 -7796 -4318
rect -7779 -4322 -7775 -4318
rect -7843 -4343 -7839 -4339
rect -7822 -4343 -7818 -4339
rect -6365 -4440 -6361 -4436
rect -6344 -4440 -6340 -4436
rect -6429 -4447 -6425 -4443
rect -6408 -4447 -6404 -4443
rect -6396 -4447 -6392 -4443
rect -6375 -4447 -6371 -4443
rect -5887 -4455 -5883 -4451
rect -5863 -4455 -5859 -4451
rect -5855 -4455 -5851 -4451
rect -5831 -4455 -5827 -4451
rect -5728 -4479 -5724 -4475
rect -5707 -4479 -5703 -4475
rect -6063 -4526 -6059 -4522
rect -6011 -4526 -6007 -4522
rect -5959 -4526 -5955 -4522
rect -5907 -4526 -5903 -4522
rect -7875 -4685 -7871 -4681
rect -7875 -4706 -7871 -4702
rect -7875 -4736 -7871 -4732
rect -7735 -4747 -7731 -4743
rect -7714 -4747 -7710 -4743
rect -7875 -4757 -7871 -4753
rect -8045 -4792 -8041 -4788
rect -8021 -4792 -8017 -4788
rect -8013 -4792 -8009 -4788
rect -7989 -4792 -7985 -4788
rect -7546 -4834 -7542 -4830
rect -7525 -4834 -7521 -4830
rect -7589 -4855 -7585 -4851
rect -7568 -4855 -7564 -4851
rect -8221 -4863 -8217 -4859
rect -8169 -4863 -8165 -4859
rect -8117 -4863 -8113 -4859
rect -8065 -4863 -8061 -4859
rect -7393 -4930 -7389 -4926
rect -7372 -4930 -7368 -4926
rect -7457 -4937 -7453 -4933
rect -7436 -4937 -7432 -4933
rect -7424 -4937 -7420 -4933
rect -7403 -4937 -7399 -4933
rect -7545 -5039 -7541 -5035
rect -7524 -5039 -7520 -5035
rect -7247 -5043 -7243 -5039
rect -7226 -5043 -7222 -5039
rect -7311 -5050 -7307 -5046
rect -7290 -5050 -7286 -5046
rect -7278 -5050 -7274 -5046
rect -7257 -5050 -7253 -5046
rect -7588 -5060 -7584 -5056
rect -7567 -5060 -7563 -5056
rect -8032 -5104 -8028 -5100
rect -8008 -5104 -8004 -5100
rect -8000 -5104 -7996 -5100
rect -7976 -5104 -7972 -5100
rect -6806 -5064 -6802 -5060
rect -6782 -5064 -6778 -5060
rect -6774 -5064 -6770 -5060
rect -6750 -5064 -6746 -5060
rect -6694 -5099 -6690 -5095
rect -6673 -5099 -6669 -5095
rect -6982 -5135 -6978 -5131
rect -6930 -5135 -6926 -5131
rect -6878 -5135 -6874 -5131
rect -6826 -5135 -6822 -5131
rect -8208 -5175 -8204 -5171
rect -8156 -5175 -8152 -5171
rect -8104 -5175 -8100 -5171
rect -8052 -5175 -8048 -5171
rect -7806 -5171 -7802 -5167
rect -7785 -5171 -7781 -5167
rect -7849 -5192 -7845 -5188
rect -7828 -5192 -7824 -5188
rect -7897 -5447 -7893 -5443
rect -7897 -5468 -7893 -5464
rect -8045 -5498 -8041 -5494
rect -8021 -5498 -8017 -5494
rect -8013 -5498 -8009 -5494
rect -7989 -5498 -7985 -5494
rect -7897 -5498 -7893 -5494
rect -7757 -5509 -7753 -5505
rect -7736 -5509 -7732 -5505
rect -7897 -5519 -7893 -5515
rect -8221 -5569 -8217 -5565
rect -8169 -5569 -8165 -5565
rect -8117 -5569 -8113 -5565
rect -8065 -5569 -8061 -5565
rect -7634 -5614 -7630 -5610
rect -7613 -5614 -7609 -5610
rect -7677 -5635 -7673 -5631
rect -7656 -5635 -7652 -5631
rect -8042 -5747 -8038 -5743
rect -8018 -5747 -8014 -5743
rect -8010 -5747 -8006 -5743
rect -7986 -5747 -7982 -5743
rect -6990 -5718 -6986 -5714
rect -6966 -5718 -6962 -5714
rect -6958 -5718 -6954 -5714
rect -6934 -5718 -6930 -5714
rect -7499 -5773 -7495 -5769
rect -7478 -5773 -7474 -5769
rect -7563 -5780 -7559 -5776
rect -7542 -5780 -7538 -5776
rect -7530 -5780 -7526 -5776
rect -7509 -5780 -7505 -5776
rect -6830 -5774 -6826 -5770
rect -6809 -5774 -6805 -5770
rect -7166 -5789 -7162 -5785
rect -7114 -5789 -7110 -5785
rect -7062 -5789 -7058 -5785
rect -7010 -5789 -7006 -5785
rect -7803 -5794 -7799 -5790
rect -7782 -5794 -7778 -5790
rect -8218 -5818 -8214 -5814
rect -8166 -5818 -8162 -5814
rect -8114 -5818 -8110 -5814
rect -8062 -5818 -8058 -5814
rect -7846 -5815 -7842 -5811
rect -7825 -5815 -7821 -5811
rect -7267 -5958 -7263 -5954
rect -7243 -5958 -7239 -5954
rect -7235 -5958 -7231 -5954
rect -7211 -5958 -7207 -5954
rect -7131 -5996 -7127 -5992
rect -7110 -5996 -7106 -5992
rect -7443 -6029 -7439 -6025
rect -7391 -6029 -7387 -6025
rect -7339 -6029 -7335 -6025
rect -7287 -6029 -7283 -6025
rect -7667 -6058 -7663 -6054
rect -7643 -6058 -7639 -6054
rect -7635 -6058 -7631 -6054
rect -7611 -6058 -7607 -6054
rect -7843 -6129 -7839 -6125
rect -7791 -6129 -7787 -6125
rect -7739 -6129 -7735 -6125
rect -7687 -6129 -7683 -6125
rect -7555 -6241 -7551 -6237
rect -7534 -6241 -7530 -6237
<< nsubstratencontact >>
rect -2923 -483 -2919 -479
rect -2906 -483 -2902 -479
rect -2896 -483 -2892 -479
rect -2879 -483 -2875 -479
rect -2861 -553 -2857 -549
rect -2844 -553 -2840 -549
rect -2503 -595 -2499 -591
rect -2447 -582 -2443 -578
rect -2430 -582 -2426 -578
rect -2503 -612 -2499 -608
rect -2503 -646 -2499 -642
rect -2293 -644 -2289 -640
rect -2276 -644 -2272 -640
rect -1796 -652 -1792 -648
rect -1774 -652 -1770 -648
rect -1764 -652 -1760 -648
rect -1742 -652 -1738 -648
rect -2503 -663 -2499 -659
rect -1997 -660 -1993 -656
rect -1975 -660 -1971 -656
rect -1945 -660 -1941 -656
rect -1923 -660 -1919 -656
rect -1893 -660 -1889 -656
rect -1871 -660 -1867 -656
rect -1841 -660 -1837 -656
rect -1819 -660 -1815 -656
rect -2244 -692 -2240 -688
rect -2227 -692 -2223 -688
rect -8119 -2975 -8115 -2971
rect -8097 -2975 -8093 -2971
rect -8087 -2975 -8083 -2971
rect -8065 -2975 -8061 -2971
rect -8320 -2983 -8316 -2979
rect -8298 -2983 -8294 -2979
rect -8268 -2983 -8264 -2979
rect -8246 -2983 -8242 -2979
rect -8216 -2983 -8212 -2979
rect -8194 -2983 -8190 -2979
rect -8164 -2983 -8160 -2979
rect -8142 -2983 -8138 -2979
rect -7795 -3068 -7791 -3064
rect -7739 -3055 -7735 -3051
rect -7722 -3055 -7718 -3051
rect -7795 -3085 -7791 -3081
rect -7635 -3080 -7631 -3076
rect -7618 -3080 -7614 -3076
rect -7608 -3080 -7604 -3076
rect -7591 -3080 -7587 -3076
rect -7795 -3119 -7791 -3115
rect -7490 -3118 -7486 -3114
rect -7473 -3118 -7469 -3114
rect -7463 -3118 -7459 -3114
rect -7446 -3118 -7442 -3114
rect -7795 -3136 -7791 -3132
rect -7297 -3134 -7293 -3130
rect -7280 -3134 -7276 -3130
rect -7270 -3134 -7266 -3130
rect -7253 -3134 -7249 -3130
rect -7151 -3132 -7147 -3128
rect -7134 -3132 -7130 -3128
rect -7124 -3132 -7120 -3128
rect -7107 -3132 -7103 -3128
rect -7007 -3136 -7003 -3132
rect -6990 -3136 -6986 -3132
rect -6980 -3136 -6976 -3132
rect -6963 -3136 -6959 -3132
rect -6852 -3138 -6848 -3134
rect -6835 -3138 -6831 -3134
rect -6825 -3138 -6821 -3134
rect -6808 -3138 -6804 -3134
rect -7573 -3150 -7569 -3146
rect -7556 -3150 -7552 -3146
rect -6717 -3146 -6713 -3142
rect -6700 -3146 -6696 -3142
rect -6690 -3146 -6686 -3142
rect -6673 -3146 -6669 -3142
rect -7428 -3188 -7424 -3184
rect -7411 -3188 -7407 -3184
rect -7853 -3241 -7849 -3237
rect -7836 -3241 -7832 -3237
rect -7826 -3241 -7822 -3237
rect -7809 -3241 -7805 -3237
rect -7235 -3204 -7231 -3200
rect -7218 -3204 -7214 -3200
rect -7089 -3202 -7085 -3198
rect -7072 -3202 -7068 -3198
rect -6945 -3206 -6941 -3202
rect -6928 -3206 -6924 -3202
rect -8105 -3279 -8101 -3275
rect -8083 -3279 -8079 -3275
rect -8073 -3279 -8069 -3275
rect -8051 -3279 -8047 -3275
rect -8306 -3287 -8302 -3283
rect -8284 -3287 -8280 -3283
rect -8254 -3287 -8250 -3283
rect -8232 -3287 -8228 -3283
rect -8202 -3287 -8198 -3283
rect -8180 -3287 -8176 -3283
rect -8150 -3287 -8146 -3283
rect -8128 -3287 -8124 -3283
rect -6790 -3208 -6786 -3204
rect -6773 -3208 -6769 -3204
rect -6556 -3202 -6552 -3198
rect -6539 -3202 -6535 -3198
rect -6655 -3216 -6651 -3212
rect -6638 -3216 -6634 -3212
rect -7791 -3311 -7787 -3307
rect -7774 -3311 -7770 -3307
rect -6507 -3250 -6503 -3246
rect -6490 -3250 -6486 -3246
rect -6394 -3258 -6390 -3254
rect -6377 -3258 -6373 -3254
rect -6345 -3306 -6341 -3302
rect -6328 -3306 -6324 -3302
rect -6236 -3314 -6232 -3310
rect -6219 -3314 -6215 -3310
rect -6187 -3362 -6183 -3358
rect -6170 -3362 -6166 -3358
rect -6070 -3390 -6066 -3386
rect -6053 -3390 -6049 -3386
rect -5719 -3429 -5715 -3425
rect -5697 -3429 -5693 -3425
rect -5687 -3429 -5683 -3425
rect -5665 -3429 -5661 -3425
rect -6021 -3438 -6017 -3434
rect -6004 -3438 -6000 -3434
rect -5920 -3437 -5916 -3433
rect -5898 -3437 -5894 -3433
rect -5868 -3437 -5864 -3433
rect -5846 -3437 -5842 -3433
rect -5816 -3437 -5812 -3433
rect -5794 -3437 -5790 -3433
rect -5764 -3437 -5760 -3433
rect -5742 -3437 -5738 -3433
rect -5550 -3471 -5546 -3467
rect -5533 -3471 -5529 -3467
rect -8050 -3887 -8046 -3883
rect -8028 -3887 -8024 -3883
rect -8018 -3887 -8014 -3883
rect -7996 -3887 -7992 -3883
rect -8251 -3895 -8247 -3891
rect -8229 -3895 -8225 -3891
rect -8199 -3895 -8195 -3891
rect -8177 -3895 -8173 -3891
rect -8147 -3895 -8143 -3891
rect -8125 -3895 -8121 -3891
rect -8095 -3895 -8091 -3891
rect -8073 -3895 -8069 -3891
rect -7627 -3895 -7623 -3891
rect -7610 -3895 -7606 -3891
rect -7600 -3895 -7596 -3891
rect -7583 -3895 -7579 -3891
rect -7458 -3894 -7454 -3890
rect -7441 -3894 -7437 -3890
rect -7431 -3894 -7427 -3890
rect -7414 -3894 -7410 -3890
rect -7294 -3892 -7290 -3888
rect -7277 -3892 -7273 -3888
rect -7267 -3892 -7263 -3888
rect -7250 -3892 -7246 -3888
rect -7154 -3894 -7150 -3890
rect -7137 -3894 -7133 -3890
rect -7127 -3894 -7123 -3890
rect -7110 -3894 -7106 -3890
rect -7789 -3919 -7785 -3915
rect -7733 -3906 -7729 -3902
rect -7716 -3906 -7712 -3902
rect -7003 -3907 -6999 -3903
rect -6986 -3907 -6982 -3903
rect -6976 -3907 -6972 -3903
rect -6959 -3907 -6955 -3903
rect -7789 -3936 -7785 -3932
rect -7789 -3970 -7785 -3966
rect -7565 -3965 -7561 -3961
rect -7548 -3965 -7544 -3961
rect -7396 -3964 -7392 -3960
rect -7379 -3964 -7375 -3960
rect -7232 -3962 -7228 -3958
rect -7215 -3962 -7211 -3958
rect -6693 -3949 -6689 -3945
rect -6676 -3949 -6672 -3945
rect -7092 -3964 -7088 -3960
rect -7075 -3964 -7071 -3960
rect -7789 -3987 -7785 -3983
rect -6941 -3977 -6937 -3973
rect -6924 -3977 -6920 -3973
rect -6644 -3997 -6640 -3993
rect -6627 -3997 -6623 -3993
rect -6840 -4111 -6836 -4107
rect -6823 -4111 -6819 -4107
rect -6813 -4111 -6809 -4107
rect -6796 -4111 -6792 -4107
rect -8033 -4128 -8029 -4124
rect -8011 -4128 -8007 -4124
rect -8001 -4128 -7997 -4124
rect -7979 -4128 -7975 -4124
rect -8234 -4136 -8230 -4132
rect -8212 -4136 -8208 -4132
rect -8182 -4136 -8178 -4132
rect -8160 -4136 -8156 -4132
rect -8130 -4136 -8126 -4132
rect -8108 -4136 -8104 -4132
rect -8078 -4136 -8074 -4132
rect -8056 -4136 -8052 -4132
rect -7860 -4156 -7856 -4152
rect -7843 -4156 -7839 -4152
rect -7833 -4156 -7829 -4152
rect -7816 -4156 -7812 -4152
rect -6559 -4159 -6555 -4155
rect -6542 -4159 -6538 -4155
rect -6778 -4181 -6774 -4177
rect -6761 -4181 -6757 -4177
rect -7798 -4226 -7794 -4222
rect -7781 -4226 -7777 -4222
rect -6510 -4207 -6506 -4203
rect -6493 -4207 -6489 -4203
rect -6412 -4319 -6408 -4315
rect -6395 -4319 -6391 -4315
rect -6363 -4367 -6359 -4363
rect -6346 -4367 -6342 -4363
rect -5886 -4354 -5882 -4350
rect -5864 -4354 -5860 -4350
rect -5854 -4354 -5850 -4350
rect -5832 -4354 -5828 -4350
rect -6087 -4362 -6083 -4358
rect -6065 -4362 -6061 -4358
rect -6035 -4362 -6031 -4358
rect -6013 -4362 -6009 -4358
rect -5983 -4362 -5979 -4358
rect -5961 -4362 -5957 -4358
rect -5931 -4362 -5927 -4358
rect -5909 -4362 -5905 -4358
rect -5726 -4383 -5722 -4379
rect -5709 -4383 -5705 -4379
rect -7606 -4668 -7602 -4664
rect -7589 -4668 -7585 -4664
rect -7579 -4668 -7575 -4664
rect -7562 -4668 -7558 -4664
rect -7789 -4687 -7785 -4683
rect -8044 -4691 -8040 -4687
rect -8022 -4691 -8018 -4687
rect -8012 -4691 -8008 -4687
rect -7990 -4691 -7986 -4687
rect -8245 -4699 -8241 -4695
rect -8223 -4699 -8219 -4695
rect -8193 -4699 -8189 -4695
rect -8171 -4699 -8167 -4695
rect -8141 -4699 -8137 -4695
rect -8119 -4699 -8115 -4695
rect -8089 -4699 -8085 -4695
rect -8067 -4699 -8063 -4695
rect -7733 -4674 -7729 -4670
rect -7716 -4674 -7712 -4670
rect -7789 -4704 -7785 -4700
rect -7789 -4738 -7785 -4734
rect -7544 -4738 -7540 -4734
rect -7527 -4738 -7523 -4734
rect -7789 -4755 -7785 -4751
rect -7440 -4809 -7436 -4805
rect -7423 -4809 -7419 -4805
rect -7605 -4873 -7601 -4869
rect -7588 -4873 -7584 -4869
rect -7578 -4873 -7574 -4869
rect -7561 -4873 -7557 -4869
rect -7391 -4857 -7387 -4853
rect -7374 -4857 -7370 -4853
rect -7294 -4922 -7290 -4918
rect -7277 -4922 -7273 -4918
rect -7543 -4943 -7539 -4939
rect -7526 -4943 -7522 -4939
rect -8031 -5003 -8027 -4999
rect -8009 -5003 -8005 -4999
rect -7999 -5003 -7995 -4999
rect -7977 -5003 -7973 -4999
rect -7866 -5005 -7862 -5001
rect -7849 -5005 -7845 -5001
rect -7839 -5005 -7835 -5001
rect -7822 -5005 -7818 -5001
rect -8232 -5011 -8228 -5007
rect -8210 -5011 -8206 -5007
rect -8180 -5011 -8176 -5007
rect -8158 -5011 -8154 -5007
rect -8128 -5011 -8124 -5007
rect -8106 -5011 -8102 -5007
rect -8076 -5011 -8072 -5007
rect -8054 -5011 -8050 -5007
rect -7245 -4970 -7241 -4966
rect -7228 -4970 -7224 -4966
rect -6805 -4963 -6801 -4959
rect -6783 -4963 -6779 -4959
rect -6773 -4963 -6769 -4959
rect -6751 -4963 -6747 -4959
rect -7006 -4971 -7002 -4967
rect -6984 -4971 -6980 -4967
rect -6954 -4971 -6950 -4967
rect -6932 -4971 -6928 -4967
rect -6902 -4971 -6898 -4967
rect -6880 -4971 -6876 -4967
rect -6850 -4971 -6846 -4967
rect -6828 -4971 -6824 -4967
rect -6692 -5003 -6688 -4999
rect -6675 -5003 -6671 -4999
rect -7804 -5075 -7800 -5071
rect -7787 -5075 -7783 -5071
rect -8044 -5397 -8040 -5393
rect -8022 -5397 -8018 -5393
rect -8012 -5397 -8008 -5393
rect -7990 -5397 -7986 -5393
rect -8245 -5405 -8241 -5401
rect -8223 -5405 -8219 -5401
rect -8193 -5405 -8189 -5401
rect -8171 -5405 -8167 -5401
rect -8141 -5405 -8137 -5401
rect -8119 -5405 -8115 -5401
rect -8089 -5405 -8085 -5401
rect -8067 -5405 -8063 -5401
rect -7811 -5449 -7807 -5445
rect -7755 -5436 -7751 -5432
rect -7738 -5436 -7734 -5432
rect -7811 -5466 -7807 -5462
rect -7694 -5448 -7690 -5444
rect -7677 -5448 -7673 -5444
rect -7667 -5448 -7663 -5444
rect -7650 -5448 -7646 -5444
rect -7811 -5500 -7807 -5496
rect -7811 -5517 -7807 -5513
rect -7632 -5518 -7628 -5514
rect -7615 -5518 -7611 -5514
rect -6989 -5617 -6985 -5613
rect -6967 -5617 -6963 -5613
rect -6957 -5617 -6953 -5613
rect -6935 -5617 -6931 -5613
rect -7863 -5628 -7859 -5624
rect -7846 -5628 -7842 -5624
rect -7836 -5628 -7832 -5624
rect -7819 -5628 -7815 -5624
rect -7190 -5625 -7186 -5621
rect -7168 -5625 -7164 -5621
rect -7138 -5625 -7134 -5621
rect -7116 -5625 -7112 -5621
rect -7086 -5625 -7082 -5621
rect -7064 -5625 -7060 -5621
rect -7034 -5625 -7030 -5621
rect -7012 -5625 -7008 -5621
rect -8041 -5646 -8037 -5642
rect -8019 -5646 -8015 -5642
rect -8009 -5646 -8005 -5642
rect -7987 -5646 -7983 -5642
rect -8242 -5654 -8238 -5650
rect -8220 -5654 -8216 -5650
rect -8190 -5654 -8186 -5650
rect -8168 -5654 -8164 -5650
rect -8138 -5654 -8134 -5650
rect -8116 -5654 -8112 -5650
rect -8086 -5654 -8082 -5650
rect -8064 -5654 -8060 -5650
rect -7546 -5652 -7542 -5648
rect -7529 -5652 -7525 -5648
rect -7801 -5698 -7797 -5694
rect -7784 -5698 -7780 -5694
rect -7497 -5700 -7493 -5696
rect -7480 -5700 -7476 -5696
rect -6828 -5678 -6824 -5674
rect -6811 -5678 -6807 -5674
rect -7266 -5857 -7262 -5853
rect -7244 -5857 -7240 -5853
rect -7234 -5857 -7230 -5853
rect -7212 -5857 -7208 -5853
rect -7467 -5865 -7463 -5861
rect -7445 -5865 -7441 -5861
rect -7415 -5865 -7411 -5861
rect -7393 -5865 -7389 -5861
rect -7363 -5865 -7359 -5861
rect -7341 -5865 -7337 -5861
rect -7311 -5865 -7307 -5861
rect -7289 -5865 -7285 -5861
rect -7129 -5900 -7125 -5896
rect -7112 -5900 -7108 -5896
rect -7666 -5957 -7662 -5953
rect -7644 -5957 -7640 -5953
rect -7634 -5957 -7630 -5953
rect -7612 -5957 -7608 -5953
rect -7867 -5965 -7863 -5961
rect -7845 -5965 -7841 -5961
rect -7815 -5965 -7811 -5961
rect -7793 -5965 -7789 -5961
rect -7763 -5965 -7759 -5961
rect -7741 -5965 -7737 -5961
rect -7711 -5965 -7707 -5961
rect -7689 -5965 -7685 -5961
rect -7553 -6145 -7549 -6141
rect -7536 -6145 -7532 -6141
<< polysilicon >>
rect -2913 -510 -2911 -506
rect -2886 -510 -2884 -506
rect -2913 -555 -2911 -530
rect -2886 -546 -2884 -530
rect -2894 -584 -2892 -557
rect -2851 -560 -2849 -557
rect -2555 -580 -2471 -578
rect -2894 -608 -2892 -604
rect -2851 -627 -2849 -600
rect -2581 -603 -2578 -601
rect -2568 -603 -2540 -601
rect -2520 -603 -2515 -601
rect -2473 -605 -2471 -580
rect -2437 -592 -2435 -586
rect -2473 -618 -2471 -615
rect -2555 -625 -2471 -623
rect -2894 -639 -2892 -630
rect -2473 -638 -2471 -625
rect -2437 -630 -2435 -612
rect -2851 -641 -2849 -638
rect -2437 -647 -2435 -640
rect -2473 -651 -2471 -648
rect -2581 -654 -2578 -652
rect -2568 -654 -2540 -652
rect -2520 -654 -2515 -652
rect -2283 -658 -2281 -648
rect -2894 -662 -2892 -659
rect -1784 -660 -1782 -656
rect -1752 -660 -1750 -656
rect -1985 -668 -1983 -664
rect -1933 -668 -1931 -664
rect -1881 -668 -1879 -664
rect -1829 -668 -1827 -664
rect -2283 -684 -2281 -678
rect -2283 -686 -2263 -684
rect -2283 -706 -2281 -697
rect -2283 -731 -2281 -725
rect -2298 -733 -2281 -731
rect -2298 -750 -2296 -733
rect -2265 -750 -2263 -686
rect -2234 -702 -2232 -696
rect -1985 -717 -1983 -708
rect -1933 -717 -1931 -708
rect -1881 -717 -1879 -708
rect -1829 -717 -1827 -708
rect -1784 -720 -1782 -700
rect -1752 -720 -1750 -700
rect -2234 -740 -2232 -722
rect -1985 -730 -1983 -726
rect -1933 -730 -1931 -726
rect -2234 -757 -2232 -750
rect -2298 -764 -2296 -760
rect -2265 -764 -2263 -760
rect -1881 -744 -1879 -735
rect -1829 -744 -1827 -735
rect -1784 -744 -1782 -740
rect -1752 -744 -1750 -740
rect -1881 -767 -1879 -764
rect -1829 -767 -1827 -764
rect -1985 -779 -1983 -770
rect -1933 -779 -1931 -770
rect -1985 -791 -1983 -783
rect -1933 -791 -1931 -783
rect -1881 -791 -1879 -783
rect -1829 -791 -1827 -783
rect -1985 -815 -1983 -811
rect -1933 -815 -1931 -811
rect -1881 -815 -1879 -811
rect -1829 -815 -1827 -811
rect -8107 -2983 -8105 -2979
rect -8075 -2983 -8073 -2979
rect -8308 -2991 -8306 -2987
rect -8256 -2991 -8254 -2987
rect -8204 -2991 -8202 -2987
rect -8152 -2991 -8150 -2987
rect -8308 -3040 -8306 -3031
rect -8256 -3040 -8254 -3031
rect -8204 -3040 -8202 -3031
rect -8152 -3040 -8150 -3031
rect -8107 -3043 -8105 -3023
rect -8075 -3043 -8073 -3023
rect -8308 -3053 -8306 -3049
rect -8256 -3053 -8254 -3049
rect -8204 -3067 -8202 -3058
rect -8152 -3067 -8150 -3058
rect -7847 -3053 -7763 -3051
rect -8107 -3067 -8105 -3063
rect -8075 -3067 -8073 -3063
rect -7873 -3076 -7870 -3074
rect -7860 -3076 -7832 -3074
rect -7812 -3076 -7807 -3074
rect -7765 -3080 -7763 -3053
rect -7729 -3065 -7727 -3059
rect -8204 -3090 -8202 -3087
rect -8152 -3090 -8150 -3087
rect -7765 -3091 -7763 -3088
rect -8308 -3102 -8306 -3093
rect -8256 -3102 -8254 -3093
rect -7847 -3098 -7763 -3096
rect -8308 -3114 -8306 -3106
rect -8256 -3114 -8254 -3106
rect -8204 -3114 -8202 -3106
rect -8152 -3114 -8150 -3106
rect -7765 -3111 -7763 -3098
rect -7729 -3103 -7727 -3085
rect -7625 -3107 -7623 -3103
rect -7598 -3107 -7596 -3103
rect -7729 -3120 -7727 -3113
rect -7765 -3124 -7763 -3121
rect -7873 -3127 -7870 -3125
rect -7860 -3127 -7832 -3125
rect -7812 -3127 -7807 -3125
rect -8308 -3138 -8306 -3134
rect -8256 -3138 -8254 -3134
rect -8204 -3138 -8202 -3134
rect -8152 -3138 -8150 -3134
rect -7625 -3152 -7623 -3127
rect -7598 -3143 -7596 -3127
rect -7480 -3145 -7478 -3141
rect -7453 -3145 -7451 -3141
rect -7606 -3181 -7604 -3154
rect -7563 -3157 -7561 -3154
rect -7287 -3161 -7285 -3157
rect -7260 -3161 -7258 -3157
rect -7141 -3159 -7139 -3155
rect -7114 -3159 -7112 -3155
rect -7480 -3190 -7478 -3165
rect -7453 -3181 -7451 -3165
rect -6997 -3163 -6995 -3159
rect -6970 -3163 -6968 -3159
rect -7606 -3205 -7604 -3201
rect -7563 -3224 -7561 -3197
rect -7461 -3219 -7459 -3192
rect -7418 -3195 -7416 -3192
rect -7606 -3236 -7604 -3227
rect -7563 -3238 -7561 -3235
rect -7287 -3206 -7285 -3181
rect -7260 -3197 -7258 -3181
rect -7141 -3204 -7139 -3179
rect -7114 -3195 -7112 -3179
rect -6842 -3165 -6840 -3161
rect -6815 -3165 -6813 -3161
rect -7268 -3235 -7266 -3208
rect -7225 -3211 -7223 -3208
rect -7461 -3243 -7459 -3239
rect -7606 -3259 -7604 -3256
rect -7418 -3262 -7416 -3235
rect -7122 -3233 -7120 -3206
rect -7079 -3209 -7077 -3206
rect -6997 -3208 -6995 -3183
rect -6970 -3199 -6968 -3183
rect -6707 -3173 -6705 -3169
rect -6680 -3173 -6678 -3169
rect -7268 -3259 -7266 -3255
rect -7843 -3268 -7841 -3264
rect -7816 -3268 -7814 -3264
rect -8093 -3287 -8091 -3283
rect -8061 -3287 -8059 -3283
rect -8294 -3295 -8292 -3291
rect -8242 -3295 -8240 -3291
rect -8190 -3295 -8188 -3291
rect -8138 -3295 -8136 -3291
rect -7461 -3274 -7459 -3265
rect -7843 -3313 -7841 -3288
rect -7816 -3304 -7814 -3288
rect -7418 -3276 -7416 -3273
rect -7225 -3278 -7223 -3251
rect -6842 -3210 -6840 -3185
rect -6815 -3201 -6813 -3185
rect -6978 -3237 -6976 -3210
rect -6935 -3213 -6933 -3210
rect -7122 -3257 -7120 -3253
rect -7079 -3276 -7077 -3249
rect -6823 -3239 -6821 -3212
rect -6780 -3215 -6778 -3212
rect -6978 -3261 -6976 -3257
rect -7268 -3290 -7266 -3281
rect -7122 -3288 -7120 -3279
rect -6935 -3280 -6933 -3253
rect -6707 -3218 -6705 -3193
rect -6680 -3209 -6678 -3193
rect -6546 -3216 -6544 -3206
rect -6688 -3247 -6686 -3220
rect -6645 -3223 -6643 -3220
rect -6823 -3263 -6821 -3259
rect -7461 -3297 -7459 -3294
rect -7225 -3292 -7223 -3289
rect -7079 -3290 -7077 -3287
rect -6978 -3292 -6976 -3283
rect -6780 -3282 -6778 -3255
rect -6546 -3242 -6544 -3236
rect -6546 -3244 -6526 -3242
rect -6688 -3271 -6686 -3267
rect -7268 -3313 -7266 -3310
rect -7122 -3311 -7120 -3308
rect -6935 -3294 -6933 -3291
rect -6823 -3294 -6821 -3285
rect -6645 -3290 -6643 -3263
rect -6546 -3264 -6544 -3255
rect -6546 -3289 -6544 -3283
rect -6978 -3315 -6976 -3312
rect -6780 -3296 -6778 -3293
rect -6688 -3302 -6686 -3293
rect -6561 -3291 -6544 -3289
rect -8294 -3344 -8292 -3335
rect -8242 -3344 -8240 -3335
rect -8190 -3344 -8188 -3335
rect -8138 -3344 -8136 -3335
rect -8093 -3347 -8091 -3327
rect -8061 -3347 -8059 -3327
rect -7824 -3342 -7822 -3315
rect -7781 -3318 -7779 -3315
rect -8294 -3357 -8292 -3353
rect -8242 -3357 -8240 -3353
rect -8190 -3371 -8188 -3362
rect -8138 -3371 -8136 -3362
rect -6823 -3317 -6821 -3314
rect -6645 -3304 -6643 -3301
rect -6561 -3308 -6559 -3291
rect -6528 -3308 -6526 -3244
rect -6497 -3260 -6495 -3254
rect -6384 -3272 -6382 -3262
rect -6497 -3298 -6495 -3280
rect -6384 -3298 -6382 -3292
rect -6384 -3300 -6364 -3298
rect -6497 -3315 -6495 -3308
rect -6561 -3322 -6559 -3318
rect -6528 -3322 -6526 -3318
rect -6688 -3325 -6686 -3322
rect -6384 -3320 -6382 -3311
rect -6384 -3345 -6382 -3339
rect -6399 -3347 -6382 -3345
rect -7824 -3366 -7822 -3362
rect -8093 -3371 -8091 -3367
rect -8061 -3371 -8059 -3367
rect -7781 -3385 -7779 -3358
rect -6399 -3364 -6397 -3347
rect -6366 -3364 -6364 -3300
rect -6335 -3316 -6333 -3310
rect -6226 -3328 -6224 -3318
rect -6335 -3354 -6333 -3336
rect -6226 -3354 -6224 -3348
rect -6226 -3356 -6206 -3354
rect -6335 -3371 -6333 -3364
rect -6399 -3378 -6397 -3374
rect -6366 -3378 -6364 -3374
rect -6226 -3376 -6224 -3367
rect -8190 -3394 -8188 -3391
rect -8138 -3394 -8136 -3391
rect -7824 -3397 -7822 -3388
rect -8294 -3406 -8292 -3397
rect -8242 -3406 -8240 -3397
rect -8294 -3418 -8292 -3410
rect -8242 -3418 -8240 -3410
rect -8190 -3418 -8188 -3410
rect -8138 -3418 -8136 -3410
rect -7781 -3399 -7779 -3396
rect -6226 -3401 -6224 -3395
rect -6241 -3403 -6224 -3401
rect -7824 -3420 -7822 -3417
rect -6241 -3420 -6239 -3403
rect -6208 -3420 -6206 -3356
rect -6177 -3372 -6175 -3366
rect -6177 -3410 -6175 -3392
rect -6060 -3404 -6058 -3394
rect -6177 -3427 -6175 -3420
rect -6241 -3434 -6239 -3430
rect -6208 -3434 -6206 -3430
rect -6060 -3430 -6058 -3424
rect -6060 -3432 -6040 -3430
rect -8294 -3442 -8292 -3438
rect -8242 -3442 -8240 -3438
rect -8190 -3442 -8188 -3438
rect -8138 -3442 -8136 -3438
rect -6060 -3452 -6058 -3443
rect -6060 -3477 -6058 -3471
rect -6075 -3479 -6058 -3477
rect -6075 -3496 -6073 -3479
rect -6042 -3496 -6040 -3432
rect -5707 -3437 -5705 -3433
rect -5675 -3437 -5673 -3433
rect -6011 -3448 -6009 -3442
rect -5908 -3445 -5906 -3441
rect -5856 -3445 -5854 -3441
rect -5804 -3445 -5802 -3441
rect -5752 -3445 -5750 -3441
rect -6011 -3486 -6009 -3468
rect -5908 -3494 -5906 -3485
rect -5856 -3494 -5854 -3485
rect -5804 -3494 -5802 -3485
rect -5752 -3494 -5750 -3485
rect -6011 -3503 -6009 -3496
rect -5707 -3497 -5705 -3477
rect -5675 -3497 -5673 -3477
rect -5540 -3478 -5538 -3475
rect -6075 -3510 -6073 -3506
rect -6042 -3510 -6040 -3506
rect -5908 -3507 -5906 -3503
rect -5856 -3507 -5854 -3503
rect -5804 -3521 -5802 -3512
rect -5752 -3521 -5750 -3512
rect -5707 -3521 -5705 -3517
rect -5675 -3521 -5673 -3517
rect -5804 -3544 -5802 -3541
rect -5752 -3544 -5750 -3541
rect -5540 -3545 -5538 -3518
rect -5908 -3556 -5906 -3547
rect -5856 -3556 -5854 -3547
rect -5540 -3559 -5538 -3556
rect -5908 -3568 -5906 -3560
rect -5856 -3568 -5854 -3560
rect -5804 -3568 -5802 -3560
rect -5752 -3568 -5750 -3560
rect -5908 -3592 -5906 -3588
rect -5856 -3592 -5854 -3588
rect -5804 -3592 -5802 -3588
rect -5752 -3592 -5750 -3588
rect -8038 -3895 -8036 -3891
rect -8006 -3895 -8004 -3891
rect -8239 -3903 -8237 -3899
rect -8187 -3903 -8185 -3899
rect -8135 -3903 -8133 -3899
rect -8083 -3903 -8081 -3899
rect -7841 -3904 -7757 -3902
rect -7867 -3927 -7864 -3925
rect -7854 -3927 -7826 -3925
rect -7806 -3927 -7801 -3925
rect -7759 -3931 -7757 -3904
rect -7723 -3916 -7721 -3910
rect -8239 -3952 -8237 -3943
rect -8187 -3952 -8185 -3943
rect -8135 -3952 -8133 -3943
rect -8083 -3952 -8081 -3943
rect -8038 -3955 -8036 -3935
rect -8006 -3955 -8004 -3935
rect -7617 -3922 -7615 -3918
rect -7590 -3922 -7588 -3918
rect -7448 -3921 -7446 -3917
rect -7421 -3921 -7419 -3917
rect -7284 -3919 -7282 -3915
rect -7257 -3919 -7255 -3915
rect -7759 -3942 -7757 -3939
rect -7841 -3949 -7757 -3947
rect -8239 -3965 -8237 -3961
rect -8187 -3965 -8185 -3961
rect -8135 -3979 -8133 -3970
rect -8083 -3979 -8081 -3970
rect -7759 -3962 -7757 -3949
rect -7723 -3954 -7721 -3936
rect -7144 -3921 -7142 -3917
rect -7117 -3921 -7115 -3917
rect -8038 -3979 -8036 -3975
rect -8006 -3979 -8004 -3975
rect -7723 -3971 -7721 -3964
rect -7617 -3967 -7615 -3942
rect -7590 -3958 -7588 -3942
rect -7448 -3966 -7446 -3941
rect -7421 -3957 -7419 -3941
rect -7284 -3964 -7282 -3939
rect -7257 -3955 -7255 -3939
rect -6993 -3934 -6991 -3930
rect -6966 -3934 -6964 -3930
rect -7144 -3966 -7142 -3941
rect -7117 -3957 -7115 -3941
rect -7759 -3975 -7757 -3972
rect -7867 -3978 -7864 -3976
rect -7854 -3978 -7826 -3976
rect -7806 -3978 -7801 -3976
rect -7598 -3996 -7596 -3969
rect -7555 -3972 -7553 -3969
rect -8135 -4002 -8133 -3999
rect -8083 -4002 -8081 -3999
rect -8239 -4014 -8237 -4005
rect -8187 -4014 -8185 -4005
rect -7429 -3995 -7427 -3968
rect -7386 -3971 -7384 -3968
rect -8239 -4026 -8237 -4018
rect -8187 -4026 -8185 -4018
rect -8135 -4026 -8133 -4018
rect -8083 -4026 -8081 -4018
rect -7598 -4020 -7596 -4016
rect -7555 -4039 -7553 -4012
rect -7265 -3993 -7263 -3966
rect -7222 -3969 -7220 -3966
rect -7429 -4019 -7427 -4015
rect -7386 -4038 -7384 -4011
rect -7125 -3995 -7123 -3968
rect -7082 -3971 -7080 -3968
rect -7265 -4017 -7263 -4013
rect -7222 -4036 -7220 -4009
rect -6993 -3979 -6991 -3954
rect -6966 -3970 -6964 -3954
rect -6683 -3963 -6681 -3953
rect -6974 -4008 -6972 -3981
rect -6931 -3984 -6929 -3981
rect -7125 -4019 -7123 -4015
rect -8239 -4050 -8237 -4046
rect -8187 -4050 -8185 -4046
rect -8135 -4050 -8133 -4046
rect -8083 -4050 -8081 -4046
rect -7598 -4051 -7596 -4042
rect -7429 -4050 -7427 -4041
rect -7265 -4048 -7263 -4039
rect -7082 -4038 -7080 -4011
rect -6683 -3989 -6681 -3983
rect -6683 -3991 -6663 -3989
rect -6683 -4011 -6681 -4002
rect -6974 -4032 -6972 -4028
rect -7555 -4053 -7553 -4050
rect -7386 -4052 -7384 -4049
rect -7222 -4050 -7220 -4047
rect -7125 -4050 -7123 -4041
rect -7598 -4074 -7596 -4071
rect -7429 -4073 -7427 -4070
rect -7265 -4071 -7263 -4068
rect -7082 -4052 -7080 -4049
rect -6931 -4051 -6929 -4024
rect -6683 -4036 -6681 -4030
rect -6698 -4038 -6681 -4036
rect -6974 -4063 -6972 -4054
rect -6698 -4055 -6696 -4038
rect -6665 -4055 -6663 -3991
rect -6634 -4007 -6632 -4001
rect -6634 -4045 -6632 -4027
rect -7125 -4073 -7123 -4070
rect -6931 -4065 -6929 -4062
rect -6634 -4062 -6632 -4055
rect -6698 -4069 -6696 -4065
rect -6665 -4069 -6663 -4065
rect -6974 -4086 -6972 -4083
rect -8021 -4136 -8019 -4132
rect -7989 -4136 -7987 -4132
rect -8222 -4144 -8220 -4140
rect -8170 -4144 -8168 -4140
rect -8118 -4144 -8116 -4140
rect -8066 -4144 -8064 -4140
rect -6830 -4138 -6828 -4134
rect -6803 -4138 -6801 -4134
rect -8222 -4193 -8220 -4184
rect -8170 -4193 -8168 -4184
rect -8118 -4193 -8116 -4184
rect -8066 -4193 -8064 -4184
rect -8021 -4196 -8019 -4176
rect -7989 -4196 -7987 -4176
rect -7850 -4183 -7848 -4179
rect -7823 -4183 -7821 -4179
rect -6830 -4183 -6828 -4158
rect -6803 -4174 -6801 -4158
rect -6549 -4173 -6547 -4163
rect -8222 -4206 -8220 -4202
rect -8170 -4206 -8168 -4202
rect -8118 -4220 -8116 -4211
rect -8066 -4220 -8064 -4211
rect -8021 -4220 -8019 -4216
rect -7989 -4220 -7987 -4216
rect -7850 -4228 -7848 -4203
rect -7823 -4219 -7821 -4203
rect -6811 -4212 -6809 -4185
rect -6768 -4188 -6766 -4185
rect -8118 -4243 -8116 -4240
rect -8066 -4243 -8064 -4240
rect -8222 -4255 -8220 -4246
rect -8170 -4255 -8168 -4246
rect -7831 -4257 -7829 -4230
rect -7788 -4233 -7786 -4230
rect -6549 -4199 -6547 -4193
rect -6549 -4201 -6529 -4199
rect -6549 -4221 -6547 -4212
rect -8222 -4267 -8220 -4259
rect -8170 -4267 -8168 -4259
rect -8118 -4267 -8116 -4259
rect -8066 -4267 -8064 -4259
rect -6811 -4236 -6809 -4232
rect -6768 -4255 -6766 -4228
rect -6549 -4246 -6547 -4240
rect -6564 -4248 -6547 -4246
rect -6811 -4267 -6809 -4258
rect -6564 -4265 -6562 -4248
rect -6531 -4265 -6529 -4201
rect -6500 -4217 -6498 -4211
rect -6500 -4255 -6498 -4237
rect -7831 -4281 -7829 -4277
rect -8222 -4291 -8220 -4287
rect -8170 -4291 -8168 -4287
rect -8118 -4291 -8116 -4287
rect -8066 -4291 -8064 -4287
rect -7788 -4300 -7786 -4273
rect -6768 -4269 -6766 -4266
rect -6500 -4272 -6498 -4265
rect -6564 -4279 -6562 -4275
rect -6531 -4279 -6529 -4275
rect -6811 -4290 -6809 -4287
rect -7831 -4312 -7829 -4303
rect -7788 -4314 -7786 -4311
rect -7831 -4335 -7829 -4332
rect -6402 -4333 -6400 -4323
rect -6192 -4346 -6190 -4342
rect -6402 -4359 -6400 -4353
rect -6402 -4361 -6382 -4359
rect -6402 -4381 -6400 -4372
rect -6402 -4406 -6400 -4400
rect -6417 -4408 -6400 -4406
rect -6417 -4425 -6415 -4408
rect -6384 -4425 -6382 -4361
rect -5874 -4362 -5872 -4358
rect -5842 -4362 -5840 -4358
rect -6353 -4377 -6351 -4371
rect -6192 -4379 -6190 -4366
rect -6075 -4370 -6073 -4366
rect -6023 -4370 -6021 -4366
rect -5971 -4370 -5969 -4366
rect -5919 -4370 -5917 -4366
rect -6192 -4393 -6190 -4389
rect -6353 -4415 -6351 -4397
rect -6192 -4401 -6190 -4397
rect -6174 -4401 -6172 -4389
rect -5716 -4390 -5714 -4387
rect -6075 -4419 -6073 -4410
rect -6023 -4419 -6021 -4410
rect -5971 -4419 -5969 -4410
rect -5919 -4419 -5917 -4410
rect -6353 -4432 -6351 -4425
rect -6192 -4433 -6190 -4421
rect -6174 -4424 -6172 -4421
rect -5874 -4422 -5872 -4402
rect -5842 -4422 -5840 -4402
rect -6174 -4433 -6172 -4430
rect -6075 -4432 -6073 -4428
rect -6023 -4432 -6021 -4428
rect -6417 -4439 -6415 -4435
rect -6384 -4439 -6382 -4435
rect -6192 -4446 -6190 -4443
rect -6174 -4449 -6172 -4443
rect -5971 -4446 -5969 -4437
rect -5919 -4446 -5917 -4437
rect -5874 -4446 -5872 -4442
rect -5842 -4446 -5840 -4442
rect -5716 -4457 -5714 -4430
rect -5971 -4469 -5969 -4466
rect -5919 -4469 -5917 -4466
rect -5716 -4471 -5714 -4468
rect -6075 -4481 -6073 -4472
rect -6023 -4481 -6021 -4472
rect -6075 -4493 -6073 -4485
rect -6023 -4493 -6021 -4485
rect -5971 -4493 -5969 -4485
rect -5919 -4493 -5917 -4485
rect -6075 -4517 -6073 -4513
rect -6023 -4517 -6021 -4513
rect -5971 -4517 -5969 -4513
rect -5919 -4517 -5917 -4513
rect -7841 -4672 -7757 -4670
rect -7867 -4695 -7864 -4693
rect -7854 -4695 -7826 -4693
rect -7806 -4695 -7801 -4693
rect -8032 -4699 -8030 -4695
rect -8000 -4699 -7998 -4695
rect -8233 -4707 -8231 -4703
rect -8181 -4707 -8179 -4703
rect -8129 -4707 -8127 -4703
rect -8077 -4707 -8075 -4703
rect -7759 -4699 -7757 -4672
rect -7723 -4684 -7721 -4678
rect -7596 -4695 -7594 -4691
rect -7569 -4695 -7567 -4691
rect -7759 -4710 -7757 -4707
rect -7841 -4717 -7757 -4715
rect -7759 -4730 -7757 -4717
rect -7723 -4722 -7721 -4704
rect -8233 -4756 -8231 -4747
rect -8181 -4756 -8179 -4747
rect -8129 -4756 -8127 -4747
rect -8077 -4756 -8075 -4747
rect -8032 -4759 -8030 -4739
rect -8000 -4759 -7998 -4739
rect -7723 -4739 -7721 -4732
rect -7596 -4740 -7594 -4715
rect -7569 -4731 -7567 -4715
rect -7759 -4743 -7757 -4740
rect -7867 -4746 -7864 -4744
rect -7854 -4746 -7826 -4744
rect -7806 -4746 -7801 -4744
rect -8233 -4769 -8231 -4765
rect -8181 -4769 -8179 -4765
rect -8129 -4783 -8127 -4774
rect -8077 -4783 -8075 -4774
rect -7577 -4769 -7575 -4742
rect -7534 -4745 -7532 -4742
rect -8032 -4783 -8030 -4779
rect -8000 -4783 -7998 -4779
rect -7577 -4793 -7575 -4789
rect -8129 -4806 -8127 -4803
rect -8077 -4806 -8075 -4803
rect -8233 -4818 -8231 -4809
rect -8181 -4818 -8179 -4809
rect -7534 -4812 -7532 -4785
rect -8233 -4830 -8231 -4822
rect -8181 -4830 -8179 -4822
rect -8129 -4830 -8127 -4822
rect -8077 -4830 -8075 -4822
rect -7577 -4824 -7575 -4815
rect -7430 -4823 -7428 -4813
rect -7534 -4826 -7532 -4823
rect -7577 -4847 -7575 -4844
rect -8233 -4854 -8231 -4850
rect -8181 -4854 -8179 -4850
rect -8129 -4854 -8127 -4850
rect -8077 -4854 -8075 -4850
rect -7430 -4849 -7428 -4843
rect -7430 -4851 -7410 -4849
rect -7430 -4871 -7428 -4862
rect -7430 -4896 -7428 -4890
rect -7595 -4900 -7593 -4896
rect -7568 -4900 -7566 -4896
rect -7445 -4898 -7428 -4896
rect -7445 -4915 -7443 -4898
rect -7412 -4915 -7410 -4851
rect -7381 -4867 -7379 -4861
rect -7381 -4905 -7379 -4887
rect -7595 -4945 -7593 -4920
rect -7568 -4936 -7566 -4920
rect -7381 -4922 -7379 -4915
rect -7445 -4929 -7443 -4925
rect -7412 -4929 -7410 -4925
rect -7284 -4936 -7282 -4926
rect -7576 -4974 -7574 -4947
rect -7533 -4950 -7531 -4947
rect -7284 -4962 -7282 -4956
rect -7110 -4957 -7108 -4953
rect -7284 -4964 -7264 -4962
rect -7284 -4984 -7282 -4975
rect -7576 -4998 -7574 -4994
rect -8019 -5011 -8017 -5007
rect -7987 -5011 -7985 -5007
rect -8220 -5019 -8218 -5015
rect -8168 -5019 -8166 -5015
rect -8116 -5019 -8114 -5015
rect -8064 -5019 -8062 -5015
rect -7533 -5017 -7531 -4990
rect -7284 -5009 -7282 -5003
rect -7299 -5011 -7282 -5009
rect -7856 -5032 -7854 -5028
rect -7829 -5032 -7827 -5028
rect -7576 -5029 -7574 -5020
rect -7299 -5028 -7297 -5011
rect -7266 -5028 -7264 -4964
rect -7235 -4980 -7233 -4974
rect -6793 -4971 -6791 -4967
rect -6761 -4971 -6759 -4967
rect -7110 -4990 -7108 -4977
rect -6994 -4979 -6992 -4975
rect -6942 -4979 -6940 -4975
rect -6890 -4979 -6888 -4975
rect -6838 -4979 -6836 -4975
rect -7235 -5018 -7233 -5000
rect -7110 -5004 -7108 -5000
rect -7110 -5012 -7108 -5008
rect -7092 -5012 -7090 -5000
rect -8220 -5068 -8218 -5059
rect -8168 -5068 -8166 -5059
rect -8116 -5068 -8114 -5059
rect -8064 -5068 -8062 -5059
rect -8019 -5071 -8017 -5051
rect -7987 -5071 -7985 -5051
rect -7533 -5031 -7531 -5028
rect -7235 -5035 -7233 -5028
rect -6682 -5010 -6680 -5007
rect -6994 -5028 -6992 -5019
rect -6942 -5028 -6940 -5019
rect -6890 -5028 -6888 -5019
rect -6838 -5028 -6836 -5019
rect -6793 -5031 -6791 -5011
rect -6761 -5031 -6759 -5011
rect -7299 -5042 -7297 -5038
rect -7266 -5042 -7264 -5038
rect -7110 -5044 -7108 -5032
rect -7092 -5035 -7090 -5032
rect -6994 -5041 -6992 -5037
rect -6942 -5041 -6940 -5037
rect -7092 -5044 -7090 -5041
rect -7576 -5052 -7574 -5049
rect -8220 -5081 -8218 -5077
rect -8168 -5081 -8166 -5077
rect -8116 -5095 -8114 -5086
rect -8064 -5095 -8062 -5086
rect -7856 -5077 -7854 -5052
rect -7829 -5068 -7827 -5052
rect -7110 -5057 -7108 -5054
rect -7092 -5060 -7090 -5054
rect -8019 -5095 -8017 -5091
rect -7987 -5095 -7985 -5091
rect -7837 -5106 -7835 -5079
rect -7794 -5082 -7792 -5079
rect -6890 -5055 -6888 -5046
rect -6838 -5055 -6836 -5046
rect -6793 -5055 -6791 -5051
rect -6761 -5055 -6759 -5051
rect -6890 -5078 -6888 -5075
rect -6838 -5078 -6836 -5075
rect -6682 -5077 -6680 -5050
rect -3985 -5057 -3983 -5053
rect -8116 -5118 -8114 -5115
rect -8064 -5118 -8062 -5115
rect -8220 -5130 -8218 -5121
rect -8168 -5130 -8166 -5121
rect -6994 -5090 -6992 -5081
rect -6942 -5090 -6940 -5081
rect -6682 -5091 -6680 -5088
rect -3985 -5090 -3983 -5077
rect -6994 -5102 -6992 -5094
rect -6942 -5102 -6940 -5094
rect -6890 -5102 -6888 -5094
rect -6838 -5102 -6836 -5094
rect -3985 -5104 -3983 -5100
rect -3985 -5112 -3983 -5108
rect -3967 -5112 -3965 -5100
rect -7837 -5130 -7835 -5126
rect -8220 -5142 -8218 -5134
rect -8168 -5142 -8166 -5134
rect -8116 -5142 -8114 -5134
rect -8064 -5142 -8062 -5134
rect -7794 -5149 -7792 -5122
rect -6994 -5126 -6992 -5122
rect -6942 -5126 -6940 -5122
rect -6890 -5126 -6888 -5122
rect -6838 -5126 -6836 -5122
rect -3985 -5144 -3983 -5132
rect -3967 -5135 -3965 -5132
rect -3967 -5144 -3965 -5141
rect -7837 -5161 -7835 -5152
rect -3985 -5157 -3983 -5154
rect -3967 -5160 -3965 -5154
rect -8220 -5166 -8218 -5162
rect -8168 -5166 -8166 -5162
rect -8116 -5166 -8114 -5162
rect -8064 -5166 -8062 -5162
rect -7794 -5163 -7792 -5160
rect -7837 -5184 -7835 -5181
rect -8032 -5405 -8030 -5401
rect -8000 -5405 -7998 -5401
rect -8233 -5413 -8231 -5409
rect -8181 -5413 -8179 -5409
rect -8129 -5413 -8127 -5409
rect -8077 -5413 -8075 -5409
rect -7863 -5434 -7779 -5432
rect -8233 -5462 -8231 -5453
rect -8181 -5462 -8179 -5453
rect -8129 -5462 -8127 -5453
rect -8077 -5462 -8075 -5453
rect -8032 -5465 -8030 -5445
rect -8000 -5465 -7998 -5445
rect -7889 -5457 -7886 -5455
rect -7876 -5457 -7848 -5455
rect -7828 -5457 -7823 -5455
rect -7781 -5461 -7779 -5434
rect -7745 -5446 -7743 -5440
rect -8233 -5475 -8231 -5471
rect -8181 -5475 -8179 -5471
rect -8129 -5489 -8127 -5480
rect -8077 -5489 -8075 -5480
rect -7781 -5472 -7779 -5469
rect -7863 -5479 -7779 -5477
rect -8032 -5489 -8030 -5485
rect -8000 -5489 -7998 -5485
rect -7781 -5492 -7779 -5479
rect -7745 -5484 -7743 -5466
rect -7684 -5475 -7682 -5471
rect -7657 -5475 -7655 -5471
rect -7745 -5501 -7743 -5494
rect -7781 -5505 -7779 -5502
rect -7889 -5508 -7886 -5506
rect -7876 -5508 -7848 -5506
rect -7828 -5508 -7823 -5506
rect -8129 -5512 -8127 -5509
rect -8077 -5512 -8075 -5509
rect -8233 -5524 -8231 -5515
rect -8181 -5524 -8179 -5515
rect -7684 -5520 -7682 -5495
rect -7657 -5511 -7655 -5495
rect -8233 -5536 -8231 -5528
rect -8181 -5536 -8179 -5528
rect -8129 -5536 -8127 -5528
rect -8077 -5536 -8075 -5528
rect -7665 -5549 -7663 -5522
rect -7622 -5525 -7620 -5522
rect -8233 -5560 -8231 -5556
rect -8181 -5560 -8179 -5556
rect -8129 -5560 -8127 -5556
rect -8077 -5560 -8075 -5556
rect -7665 -5573 -7663 -5569
rect -7622 -5592 -7620 -5565
rect -7665 -5604 -7663 -5595
rect -7622 -5606 -7620 -5603
rect -7665 -5627 -7663 -5624
rect -6977 -5625 -6975 -5621
rect -6945 -5625 -6943 -5621
rect -7178 -5633 -7176 -5629
rect -7126 -5633 -7124 -5629
rect -7074 -5633 -7072 -5629
rect -7022 -5633 -7020 -5629
rect -8029 -5654 -8027 -5650
rect -7997 -5654 -7995 -5650
rect -8230 -5662 -8228 -5658
rect -8178 -5662 -8176 -5658
rect -8126 -5662 -8124 -5658
rect -8074 -5662 -8072 -5658
rect -7853 -5655 -7851 -5651
rect -7826 -5655 -7824 -5651
rect -7536 -5666 -7534 -5656
rect -8230 -5711 -8228 -5702
rect -8178 -5711 -8176 -5702
rect -8126 -5711 -8124 -5702
rect -8074 -5711 -8072 -5702
rect -8029 -5714 -8027 -5694
rect -7997 -5714 -7995 -5694
rect -7853 -5700 -7851 -5675
rect -7826 -5691 -7824 -5675
rect -7302 -5681 -7300 -5677
rect -7536 -5692 -7534 -5686
rect -7536 -5694 -7516 -5692
rect -8230 -5724 -8228 -5720
rect -8178 -5724 -8176 -5720
rect -8126 -5738 -8124 -5729
rect -8074 -5738 -8072 -5729
rect -7834 -5729 -7832 -5702
rect -7791 -5705 -7789 -5702
rect -8029 -5738 -8027 -5734
rect -7997 -5738 -7995 -5734
rect -7536 -5714 -7534 -5705
rect -7536 -5739 -7534 -5733
rect -7551 -5741 -7534 -5739
rect -7834 -5753 -7832 -5749
rect -8126 -5761 -8124 -5758
rect -8074 -5761 -8072 -5758
rect -8230 -5773 -8228 -5764
rect -8178 -5773 -8176 -5764
rect -7791 -5772 -7789 -5745
rect -7551 -5758 -7549 -5741
rect -7518 -5758 -7516 -5694
rect -7178 -5682 -7176 -5673
rect -7126 -5682 -7124 -5673
rect -7074 -5682 -7072 -5673
rect -7022 -5682 -7020 -5673
rect -6977 -5685 -6975 -5665
rect -6945 -5685 -6943 -5665
rect -6818 -5685 -6816 -5682
rect -7178 -5695 -7176 -5691
rect -7126 -5695 -7124 -5691
rect -7487 -5710 -7485 -5704
rect -7302 -5714 -7300 -5701
rect -7302 -5728 -7300 -5724
rect -7487 -5748 -7485 -5730
rect -7302 -5736 -7300 -5732
rect -7284 -5736 -7282 -5724
rect -7074 -5709 -7072 -5700
rect -7022 -5709 -7020 -5700
rect -6977 -5709 -6975 -5705
rect -6945 -5709 -6943 -5705
rect -7074 -5732 -7072 -5729
rect -7022 -5732 -7020 -5729
rect -7178 -5744 -7176 -5735
rect -7126 -5744 -7124 -5735
rect -7178 -5756 -7176 -5748
rect -7126 -5756 -7124 -5748
rect -7074 -5756 -7072 -5748
rect -7022 -5756 -7020 -5748
rect -6818 -5752 -6816 -5725
rect -7487 -5765 -7485 -5758
rect -7302 -5768 -7300 -5756
rect -7284 -5759 -7282 -5756
rect -7284 -5768 -7282 -5765
rect -7551 -5772 -7549 -5768
rect -7518 -5772 -7516 -5768
rect -8230 -5785 -8228 -5777
rect -8178 -5785 -8176 -5777
rect -8126 -5785 -8124 -5777
rect -8074 -5785 -8072 -5777
rect -7834 -5784 -7832 -5775
rect -6818 -5766 -6816 -5763
rect -7302 -5781 -7300 -5778
rect -7791 -5786 -7789 -5783
rect -7284 -5784 -7282 -5778
rect -7178 -5780 -7176 -5776
rect -7126 -5780 -7124 -5776
rect -7074 -5780 -7072 -5776
rect -7022 -5780 -7020 -5776
rect -7630 -5797 -7628 -5793
rect -8230 -5809 -8228 -5805
rect -8178 -5809 -8176 -5805
rect -8126 -5809 -8124 -5805
rect -8074 -5809 -8072 -5805
rect -7834 -5807 -7832 -5804
rect -7630 -5830 -7628 -5817
rect -7630 -5844 -7628 -5840
rect -7630 -5852 -7628 -5848
rect -7612 -5852 -7610 -5840
rect -7254 -5865 -7252 -5861
rect -7222 -5865 -7220 -5861
rect -7630 -5884 -7628 -5872
rect -7612 -5875 -7610 -5872
rect -7455 -5873 -7453 -5869
rect -7403 -5873 -7401 -5869
rect -7351 -5873 -7349 -5869
rect -7299 -5873 -7297 -5869
rect -7612 -5884 -7610 -5881
rect -7630 -5897 -7628 -5894
rect -7612 -5900 -7610 -5894
rect -7455 -5922 -7453 -5913
rect -7403 -5922 -7401 -5913
rect -7351 -5922 -7349 -5913
rect -7299 -5922 -7297 -5913
rect -7254 -5925 -7252 -5905
rect -7222 -5925 -7220 -5905
rect -7119 -5907 -7117 -5904
rect -7455 -5935 -7453 -5931
rect -7403 -5935 -7401 -5931
rect -7654 -5965 -7652 -5961
rect -7622 -5965 -7620 -5961
rect -7855 -5973 -7853 -5969
rect -7803 -5973 -7801 -5969
rect -7751 -5973 -7749 -5969
rect -7699 -5973 -7697 -5969
rect -7351 -5949 -7349 -5940
rect -7299 -5949 -7297 -5940
rect -7254 -5949 -7252 -5945
rect -7222 -5949 -7220 -5945
rect -7351 -5972 -7349 -5969
rect -7299 -5972 -7297 -5969
rect -7119 -5974 -7117 -5947
rect -7455 -5984 -7453 -5975
rect -7403 -5984 -7401 -5975
rect -7119 -5988 -7117 -5985
rect -7455 -5996 -7453 -5988
rect -7403 -5996 -7401 -5988
rect -7351 -5996 -7349 -5988
rect -7299 -5996 -7297 -5988
rect -7855 -6022 -7853 -6013
rect -7803 -6022 -7801 -6013
rect -7751 -6022 -7749 -6013
rect -7699 -6022 -7697 -6013
rect -7654 -6025 -7652 -6005
rect -7622 -6025 -7620 -6005
rect -7455 -6020 -7453 -6016
rect -7403 -6020 -7401 -6016
rect -7351 -6020 -7349 -6016
rect -7299 -6020 -7297 -6016
rect -7855 -6035 -7853 -6031
rect -7803 -6035 -7801 -6031
rect -7751 -6049 -7749 -6040
rect -7699 -6049 -7697 -6040
rect -7654 -6049 -7652 -6045
rect -7622 -6049 -7620 -6045
rect -7751 -6072 -7749 -6069
rect -7699 -6072 -7697 -6069
rect -7855 -6084 -7853 -6075
rect -7803 -6084 -7801 -6075
rect -7855 -6096 -7853 -6088
rect -7803 -6096 -7801 -6088
rect -7751 -6096 -7749 -6088
rect -7699 -6096 -7697 -6088
rect -7855 -6120 -7853 -6116
rect -7803 -6120 -7801 -6116
rect -7751 -6120 -7749 -6116
rect -7699 -6120 -7697 -6116
rect -7543 -6152 -7541 -6149
rect -7543 -6219 -7541 -6192
rect -7543 -6233 -7541 -6230
<< polycontact >>
rect -2918 -552 -2913 -547
rect -2884 -546 -2879 -542
rect -2900 -562 -2894 -557
rect -2555 -585 -2550 -580
rect -2856 -615 -2851 -610
rect -2555 -601 -2550 -596
rect -2555 -623 -2550 -618
rect -2901 -636 -2894 -631
rect -2442 -627 -2437 -622
rect -2555 -652 -2550 -647
rect -2288 -686 -2283 -681
rect -2303 -736 -2298 -731
rect -1990 -717 -1985 -712
rect -1938 -717 -1933 -712
rect -1886 -717 -1881 -712
rect -1834 -717 -1829 -712
rect -1789 -717 -1784 -712
rect -1757 -717 -1752 -712
rect -2239 -737 -2234 -732
rect -1886 -740 -1881 -735
rect -1834 -740 -1829 -735
rect -1990 -779 -1985 -774
rect -1938 -779 -1933 -774
rect -1990 -788 -1985 -783
rect -1938 -788 -1933 -783
rect -1886 -788 -1881 -783
rect -1834 -788 -1829 -783
rect -8313 -3040 -8308 -3035
rect -8261 -3040 -8256 -3035
rect -8209 -3040 -8204 -3035
rect -8157 -3040 -8152 -3035
rect -8112 -3040 -8107 -3035
rect -8080 -3040 -8075 -3035
rect -8209 -3063 -8204 -3058
rect -8157 -3063 -8152 -3058
rect -7847 -3058 -7842 -3053
rect -7847 -3074 -7842 -3069
rect -8313 -3102 -8308 -3097
rect -8261 -3102 -8256 -3097
rect -7847 -3096 -7842 -3091
rect -8313 -3111 -8308 -3106
rect -8261 -3111 -8256 -3106
rect -8209 -3111 -8204 -3106
rect -8157 -3111 -8152 -3106
rect -7734 -3100 -7729 -3095
rect -7847 -3125 -7842 -3120
rect -7630 -3149 -7625 -3144
rect -7596 -3143 -7591 -3139
rect -7612 -3159 -7606 -3154
rect -7485 -3187 -7480 -3182
rect -7451 -3181 -7446 -3177
rect -7467 -3197 -7461 -3192
rect -7568 -3212 -7563 -3207
rect -7613 -3233 -7606 -3228
rect -7292 -3203 -7287 -3198
rect -7258 -3197 -7253 -3193
rect -7146 -3201 -7141 -3196
rect -7112 -3195 -7107 -3191
rect -7002 -3205 -6997 -3200
rect -7274 -3213 -7268 -3208
rect -7128 -3211 -7122 -3206
rect -7423 -3250 -7418 -3245
rect -6968 -3199 -6963 -3195
rect -6847 -3207 -6842 -3202
rect -7468 -3271 -7461 -3266
rect -7230 -3266 -7225 -3261
rect -7848 -3310 -7843 -3305
rect -6813 -3201 -6808 -3197
rect -6984 -3215 -6978 -3210
rect -7084 -3264 -7079 -3259
rect -6829 -3217 -6823 -3212
rect -6712 -3215 -6707 -3210
rect -6940 -3268 -6935 -3263
rect -7275 -3287 -7268 -3282
rect -7129 -3285 -7122 -3280
rect -6678 -3209 -6673 -3205
rect -6694 -3225 -6688 -3220
rect -6785 -3270 -6780 -3265
rect -7814 -3304 -7809 -3300
rect -6985 -3289 -6978 -3284
rect -6551 -3244 -6546 -3239
rect -6650 -3278 -6645 -3273
rect -6830 -3291 -6823 -3286
rect -6695 -3299 -6688 -3294
rect -6566 -3294 -6561 -3289
rect -7830 -3320 -7824 -3315
rect -8299 -3344 -8294 -3339
rect -8247 -3344 -8242 -3339
rect -8195 -3344 -8190 -3339
rect -8143 -3344 -8138 -3339
rect -8098 -3344 -8093 -3339
rect -8066 -3344 -8061 -3339
rect -8195 -3367 -8190 -3362
rect -8143 -3367 -8138 -3362
rect -6502 -3295 -6497 -3290
rect -6389 -3300 -6384 -3295
rect -6404 -3350 -6399 -3345
rect -7786 -3373 -7781 -3368
rect -6340 -3351 -6335 -3346
rect -6231 -3356 -6226 -3351
rect -7831 -3394 -7824 -3389
rect -8299 -3406 -8294 -3401
rect -8247 -3406 -8242 -3401
rect -8299 -3415 -8294 -3410
rect -8247 -3415 -8242 -3410
rect -8195 -3415 -8190 -3410
rect -8143 -3415 -8138 -3410
rect -6246 -3406 -6241 -3401
rect -6182 -3407 -6177 -3402
rect -6065 -3432 -6060 -3427
rect -6080 -3482 -6075 -3477
rect -6016 -3483 -6011 -3478
rect -5913 -3494 -5908 -3489
rect -5861 -3494 -5856 -3489
rect -5809 -3494 -5804 -3489
rect -5757 -3494 -5752 -3489
rect -5712 -3494 -5707 -3489
rect -5680 -3494 -5675 -3489
rect -5809 -3517 -5804 -3512
rect -5757 -3517 -5752 -3512
rect -5545 -3533 -5540 -3528
rect -5913 -3556 -5908 -3551
rect -5861 -3556 -5856 -3551
rect -5913 -3565 -5908 -3560
rect -5861 -3565 -5856 -3560
rect -5809 -3565 -5804 -3560
rect -5757 -3565 -5752 -3560
rect -7841 -3909 -7836 -3904
rect -7841 -3925 -7836 -3920
rect -8244 -3952 -8239 -3947
rect -8192 -3952 -8187 -3947
rect -8140 -3952 -8135 -3947
rect -8088 -3952 -8083 -3947
rect -8043 -3952 -8038 -3947
rect -8011 -3952 -8006 -3947
rect -7841 -3947 -7836 -3942
rect -8140 -3975 -8135 -3970
rect -8088 -3975 -8083 -3970
rect -7728 -3951 -7723 -3946
rect -7841 -3976 -7836 -3971
rect -7622 -3964 -7617 -3959
rect -7588 -3958 -7583 -3954
rect -7453 -3963 -7448 -3958
rect -7419 -3957 -7414 -3953
rect -7289 -3961 -7284 -3956
rect -7255 -3955 -7250 -3951
rect -7149 -3963 -7144 -3958
rect -7115 -3957 -7110 -3953
rect -7604 -3974 -7598 -3969
rect -8244 -4014 -8239 -4009
rect -8192 -4014 -8187 -4009
rect -7435 -3973 -7429 -3968
rect -7271 -3971 -7265 -3966
rect -8244 -4023 -8239 -4018
rect -8192 -4023 -8187 -4018
rect -8140 -4023 -8135 -4018
rect -8088 -4023 -8083 -4018
rect -7560 -4027 -7555 -4022
rect -7391 -4026 -7386 -4021
rect -7131 -3973 -7125 -3968
rect -7227 -4024 -7222 -4019
rect -6998 -3976 -6993 -3971
rect -6964 -3970 -6959 -3966
rect -6980 -3986 -6974 -3981
rect -7087 -4026 -7082 -4021
rect -7605 -4048 -7598 -4043
rect -7436 -4047 -7429 -4042
rect -7272 -4045 -7265 -4040
rect -6688 -3991 -6683 -3986
rect -7132 -4047 -7125 -4042
rect -6936 -4039 -6931 -4034
rect -6703 -4041 -6698 -4036
rect -6981 -4060 -6974 -4055
rect -6639 -4042 -6634 -4037
rect -8227 -4193 -8222 -4188
rect -8175 -4193 -8170 -4188
rect -8123 -4193 -8118 -4188
rect -8071 -4193 -8066 -4188
rect -8026 -4193 -8021 -4188
rect -7994 -4193 -7989 -4188
rect -6835 -4180 -6830 -4175
rect -6801 -4174 -6796 -4170
rect -8123 -4216 -8118 -4211
rect -8071 -4216 -8066 -4211
rect -6817 -4190 -6811 -4185
rect -7855 -4225 -7850 -4220
rect -7821 -4219 -7816 -4215
rect -7837 -4235 -7831 -4230
rect -8227 -4255 -8222 -4250
rect -8175 -4255 -8170 -4250
rect -6554 -4201 -6549 -4196
rect -8227 -4264 -8222 -4259
rect -8175 -4264 -8170 -4259
rect -8123 -4264 -8118 -4259
rect -8071 -4264 -8066 -4259
rect -6773 -4243 -6768 -4238
rect -6569 -4251 -6564 -4246
rect -6818 -4264 -6811 -4259
rect -6505 -4252 -6500 -4247
rect -7793 -4288 -7788 -4283
rect -7838 -4309 -7831 -4304
rect -6407 -4361 -6402 -4356
rect -6422 -4411 -6417 -4406
rect -6196 -4378 -6192 -4374
rect -6178 -4394 -6174 -4390
rect -6358 -4412 -6353 -4407
rect -6080 -4419 -6075 -4414
rect -6028 -4419 -6023 -4414
rect -5976 -4419 -5971 -4414
rect -5924 -4419 -5919 -4414
rect -5879 -4419 -5874 -4414
rect -6196 -4432 -6192 -4428
rect -5847 -4419 -5842 -4414
rect -6172 -4448 -6168 -4444
rect -5976 -4442 -5971 -4437
rect -5924 -4442 -5919 -4437
rect -5721 -4445 -5716 -4440
rect -6080 -4481 -6075 -4476
rect -6028 -4481 -6023 -4476
rect -6080 -4490 -6075 -4485
rect -6028 -4490 -6023 -4485
rect -5976 -4490 -5971 -4485
rect -5924 -4490 -5919 -4485
rect -7841 -4677 -7836 -4672
rect -7841 -4693 -7836 -4688
rect -7841 -4715 -7836 -4710
rect -7728 -4719 -7723 -4714
rect -8238 -4756 -8233 -4751
rect -8186 -4756 -8181 -4751
rect -8134 -4756 -8129 -4751
rect -8082 -4756 -8077 -4751
rect -8037 -4756 -8032 -4751
rect -8005 -4756 -8000 -4751
rect -7841 -4744 -7836 -4739
rect -7601 -4737 -7596 -4732
rect -7567 -4731 -7562 -4727
rect -7583 -4747 -7577 -4742
rect -8134 -4779 -8129 -4774
rect -8082 -4779 -8077 -4774
rect -7539 -4800 -7534 -4795
rect -8238 -4818 -8233 -4813
rect -8186 -4818 -8181 -4813
rect -7584 -4821 -7577 -4816
rect -8238 -4827 -8233 -4822
rect -8186 -4827 -8181 -4822
rect -8134 -4827 -8129 -4822
rect -8082 -4827 -8077 -4822
rect -7435 -4851 -7430 -4846
rect -7450 -4901 -7445 -4896
rect -7386 -4902 -7381 -4897
rect -7600 -4942 -7595 -4937
rect -7566 -4936 -7561 -4932
rect -7582 -4952 -7576 -4947
rect -7289 -4964 -7284 -4959
rect -7538 -5005 -7533 -5000
rect -7304 -5014 -7299 -5009
rect -7583 -5026 -7576 -5021
rect -7114 -4989 -7110 -4985
rect -7240 -5015 -7235 -5010
rect -7096 -5005 -7092 -5001
rect -8225 -5068 -8220 -5063
rect -8173 -5068 -8168 -5063
rect -8121 -5068 -8116 -5063
rect -8069 -5068 -8064 -5063
rect -8024 -5068 -8019 -5063
rect -7992 -5068 -7987 -5063
rect -6999 -5028 -6994 -5023
rect -6947 -5028 -6942 -5023
rect -6895 -5028 -6890 -5023
rect -6843 -5028 -6838 -5023
rect -6798 -5028 -6793 -5023
rect -6766 -5028 -6761 -5023
rect -7114 -5043 -7110 -5039
rect -8121 -5091 -8116 -5086
rect -8069 -5091 -8064 -5086
rect -7861 -5074 -7856 -5069
rect -7090 -5059 -7086 -5055
rect -7827 -5068 -7822 -5064
rect -7843 -5084 -7837 -5079
rect -6895 -5051 -6890 -5046
rect -6843 -5051 -6838 -5046
rect -6687 -5065 -6682 -5060
rect -8225 -5130 -8220 -5125
rect -8173 -5130 -8168 -5125
rect -6999 -5090 -6994 -5085
rect -6947 -5090 -6942 -5085
rect -3989 -5089 -3985 -5085
rect -6999 -5099 -6994 -5094
rect -6947 -5099 -6942 -5094
rect -6895 -5099 -6890 -5094
rect -6843 -5099 -6838 -5094
rect -3971 -5105 -3967 -5101
rect -8225 -5139 -8220 -5134
rect -8173 -5139 -8168 -5134
rect -8121 -5139 -8116 -5134
rect -8069 -5139 -8064 -5134
rect -7799 -5137 -7794 -5132
rect -3989 -5143 -3985 -5139
rect -7844 -5158 -7837 -5153
rect -3965 -5159 -3961 -5155
rect -7863 -5439 -7858 -5434
rect -8238 -5462 -8233 -5457
rect -8186 -5462 -8181 -5457
rect -8134 -5462 -8129 -5457
rect -8082 -5462 -8077 -5457
rect -8037 -5462 -8032 -5457
rect -8005 -5462 -8000 -5457
rect -7863 -5455 -7858 -5450
rect -8134 -5485 -8129 -5480
rect -8082 -5485 -8077 -5480
rect -7863 -5477 -7858 -5472
rect -7750 -5481 -7745 -5476
rect -7863 -5506 -7858 -5501
rect -8238 -5524 -8233 -5519
rect -8186 -5524 -8181 -5519
rect -7689 -5517 -7684 -5512
rect -7655 -5511 -7650 -5507
rect -7671 -5527 -7665 -5522
rect -8238 -5533 -8233 -5528
rect -8186 -5533 -8181 -5528
rect -8134 -5533 -8129 -5528
rect -8082 -5533 -8077 -5528
rect -7627 -5580 -7622 -5575
rect -7672 -5601 -7665 -5596
rect -8235 -5711 -8230 -5706
rect -8183 -5711 -8178 -5706
rect -8131 -5711 -8126 -5706
rect -8079 -5711 -8074 -5706
rect -8034 -5711 -8029 -5706
rect -8002 -5711 -7997 -5706
rect -7858 -5697 -7853 -5692
rect -7824 -5691 -7819 -5687
rect -7541 -5694 -7536 -5689
rect -7840 -5707 -7834 -5702
rect -8131 -5734 -8126 -5729
rect -8079 -5734 -8074 -5729
rect -7556 -5744 -7551 -5739
rect -7796 -5760 -7791 -5755
rect -8235 -5773 -8230 -5768
rect -8183 -5773 -8178 -5768
rect -7183 -5682 -7178 -5677
rect -7131 -5682 -7126 -5677
rect -7079 -5682 -7074 -5677
rect -7027 -5682 -7022 -5677
rect -6982 -5682 -6977 -5677
rect -6950 -5682 -6945 -5677
rect -7306 -5713 -7302 -5709
rect -7288 -5729 -7284 -5725
rect -7492 -5745 -7487 -5740
rect -7079 -5705 -7074 -5700
rect -7027 -5705 -7022 -5700
rect -7183 -5744 -7178 -5739
rect -7131 -5744 -7126 -5739
rect -6823 -5740 -6818 -5735
rect -7183 -5753 -7178 -5748
rect -7131 -5753 -7126 -5748
rect -7079 -5753 -7074 -5748
rect -7027 -5753 -7022 -5748
rect -7306 -5767 -7302 -5763
rect -8235 -5782 -8230 -5777
rect -8183 -5782 -8178 -5777
rect -8131 -5782 -8126 -5777
rect -8079 -5782 -8074 -5777
rect -7841 -5781 -7834 -5776
rect -7282 -5783 -7278 -5779
rect -7634 -5829 -7630 -5825
rect -7616 -5845 -7612 -5841
rect -7634 -5883 -7630 -5879
rect -7610 -5899 -7606 -5895
rect -7460 -5922 -7455 -5917
rect -7408 -5922 -7403 -5917
rect -7356 -5922 -7351 -5917
rect -7304 -5922 -7299 -5917
rect -7259 -5922 -7254 -5917
rect -7227 -5922 -7222 -5917
rect -7356 -5945 -7351 -5940
rect -7304 -5945 -7299 -5940
rect -7124 -5962 -7119 -5957
rect -7460 -5984 -7455 -5979
rect -7408 -5984 -7403 -5979
rect -7460 -5993 -7455 -5988
rect -7408 -5993 -7403 -5988
rect -7356 -5993 -7351 -5988
rect -7304 -5993 -7299 -5988
rect -7860 -6022 -7855 -6017
rect -7808 -6022 -7803 -6017
rect -7756 -6022 -7751 -6017
rect -7704 -6022 -7699 -6017
rect -7659 -6022 -7654 -6017
rect -7627 -6022 -7622 -6017
rect -7756 -6045 -7751 -6040
rect -7704 -6045 -7699 -6040
rect -7860 -6084 -7855 -6079
rect -7808 -6084 -7803 -6079
rect -7860 -6093 -7855 -6088
rect -7808 -6093 -7803 -6088
rect -7756 -6093 -7751 -6088
rect -7704 -6093 -7699 -6088
rect -7548 -6207 -7543 -6202
<< metal1 >>
rect -2926 -479 -2872 -476
rect -2926 -483 -2923 -479
rect -2919 -483 -2906 -479
rect -2902 -483 -2896 -479
rect -2892 -483 -2879 -479
rect -2875 -483 -2872 -479
rect -2926 -485 -2872 -483
rect -2918 -510 -2914 -485
rect -2883 -510 -2879 -485
rect -2931 -552 -2918 -547
rect -2910 -550 -2906 -530
rect -2891 -550 -2887 -530
rect -2879 -546 -2872 -542
rect -2931 -557 -2926 -552
rect -2910 -554 -2887 -550
rect -2877 -554 -2872 -546
rect -2864 -549 -2837 -546
rect -2864 -553 -2861 -549
rect -2857 -553 -2844 -549
rect -2840 -553 -2837 -549
rect -2931 -562 -2900 -557
rect -2931 -575 -2926 -562
rect -2939 -578 -2926 -575
rect -2891 -574 -2887 -554
rect -2864 -555 -2837 -553
rect -2856 -560 -2852 -555
rect -2891 -580 -2868 -574
rect -2891 -584 -2887 -580
rect -2899 -610 -2895 -604
rect -2874 -610 -2868 -580
rect -2450 -578 -2423 -575
rect -2581 -585 -2555 -580
rect -2450 -582 -2447 -578
rect -2443 -582 -2430 -578
rect -2426 -582 -2423 -578
rect -2450 -584 -2423 -582
rect -2848 -610 -2844 -600
rect -2590 -589 -2584 -588
rect -2590 -593 -2589 -589
rect -2585 -593 -2584 -589
rect -2590 -596 -2584 -593
rect -2555 -596 -2550 -585
rect -2505 -591 -2496 -588
rect -2505 -595 -2503 -591
rect -2499 -595 -2496 -591
rect -2505 -596 -2496 -595
rect -2590 -600 -2578 -596
rect -2590 -610 -2584 -600
rect -2520 -600 -2496 -596
rect -2442 -592 -2438 -584
rect -2555 -608 -2540 -604
rect -2505 -608 -2496 -600
rect -2470 -604 -2457 -600
rect -2470 -605 -2466 -604
rect -2899 -614 -2887 -610
rect -2926 -631 -2920 -630
rect -2926 -636 -2913 -631
rect -2907 -636 -2901 -631
rect -2891 -639 -2887 -614
rect -2874 -615 -2856 -610
rect -2848 -615 -2835 -610
rect -2590 -614 -2589 -610
rect -2585 -614 -2584 -610
rect -2590 -615 -2584 -614
rect -2848 -627 -2844 -615
rect -2555 -618 -2550 -608
rect -2505 -612 -2503 -608
rect -2499 -612 -2496 -608
rect -2505 -615 -2496 -612
rect -2478 -618 -2474 -615
rect -2526 -622 -2474 -618
rect -2526 -627 -2522 -622
rect -2585 -632 -2522 -627
rect -2856 -644 -2852 -638
rect -2590 -640 -2584 -639
rect -2590 -644 -2589 -640
rect -2585 -644 -2584 -640
rect -2864 -645 -2837 -644
rect -2864 -649 -2863 -645
rect -2859 -649 -2842 -645
rect -2838 -649 -2837 -645
rect -2864 -650 -2837 -649
rect -2590 -647 -2584 -644
rect -2555 -647 -2550 -632
rect -2470 -638 -2466 -615
rect -2463 -622 -2457 -604
rect -2434 -622 -2430 -612
rect -2463 -627 -2442 -622
rect -2434 -627 -2424 -622
rect -2434 -630 -2430 -627
rect -2505 -642 -2496 -639
rect -2505 -646 -2503 -642
rect -2499 -646 -2496 -642
rect -2505 -647 -2496 -646
rect -2590 -651 -2578 -647
rect -2899 -665 -2895 -659
rect -2590 -661 -2584 -651
rect -2520 -651 -2496 -647
rect -2555 -659 -2540 -655
rect -2505 -659 -2496 -651
rect -2590 -665 -2589 -661
rect -2585 -665 -2584 -661
rect -2907 -666 -2880 -665
rect -2590 -666 -2584 -665
rect -2907 -670 -2906 -666
rect -2902 -670 -2885 -666
rect -2881 -670 -2880 -666
rect -2907 -671 -2880 -670
rect -2555 -670 -2550 -659
rect -2505 -663 -2503 -659
rect -2499 -663 -2496 -659
rect -2505 -666 -2496 -663
rect -2296 -640 -2269 -637
rect -2478 -670 -2474 -648
rect -2442 -650 -2438 -640
rect -2296 -644 -2293 -640
rect -2289 -644 -2276 -640
rect -2272 -644 -2269 -640
rect -2296 -646 -2269 -644
rect -2450 -651 -2423 -650
rect -2450 -655 -2449 -651
rect -2445 -655 -2428 -651
rect -2424 -655 -2423 -651
rect -2450 -656 -2423 -655
rect -2555 -673 -2474 -670
rect -2288 -658 -2284 -646
rect -1799 -648 -1735 -645
rect -1799 -652 -1796 -648
rect -1792 -652 -1774 -648
rect -1770 -652 -1764 -648
rect -1760 -652 -1742 -648
rect -1738 -652 -1735 -648
rect -2000 -656 -1812 -653
rect -1799 -654 -1735 -652
rect -2000 -660 -1997 -656
rect -1993 -660 -1975 -656
rect -1971 -660 -1945 -656
rect -1941 -660 -1923 -656
rect -1919 -660 -1893 -656
rect -1889 -660 -1871 -656
rect -1867 -660 -1841 -656
rect -1837 -660 -1819 -656
rect -1815 -660 -1812 -656
rect -2000 -662 -1812 -660
rect -1789 -660 -1785 -654
rect -1757 -660 -1753 -654
rect -2305 -686 -2288 -681
rect -2280 -690 -2276 -678
rect -1990 -668 -1986 -662
rect -1938 -668 -1934 -662
rect -1886 -668 -1882 -662
rect -1834 -668 -1830 -662
rect -2288 -694 -2276 -690
rect -2247 -688 -2220 -685
rect -2247 -692 -2244 -688
rect -2240 -692 -2227 -688
rect -2223 -692 -2220 -688
rect -2247 -694 -2220 -692
rect -2288 -706 -2284 -694
rect -2239 -702 -2235 -694
rect -2312 -736 -2303 -731
rect -2280 -732 -2276 -725
rect -2231 -732 -2227 -722
rect -2013 -717 -1990 -712
rect -2280 -737 -2239 -732
rect -2231 -737 -2218 -732
rect -2280 -740 -2276 -737
rect -2231 -740 -2227 -737
rect -2295 -744 -2258 -740
rect -2295 -750 -2291 -744
rect -2262 -750 -2258 -744
rect -2239 -760 -2235 -750
rect -2303 -767 -2299 -760
rect -2270 -767 -2266 -760
rect -2247 -761 -2220 -760
rect -2247 -765 -2246 -761
rect -2242 -765 -2225 -761
rect -2221 -765 -2220 -761
rect -2247 -766 -2220 -765
rect -2311 -768 -2284 -767
rect -2311 -772 -2310 -768
rect -2306 -772 -2289 -768
rect -2285 -772 -2284 -768
rect -2311 -773 -2284 -772
rect -2278 -768 -2251 -767
rect -2278 -772 -2277 -768
rect -2273 -772 -2256 -768
rect -2252 -772 -2251 -768
rect -2278 -773 -2251 -772
rect -2013 -783 -2008 -717
rect -1982 -721 -1978 -708
rect -1990 -725 -1978 -721
rect -1960 -717 -1938 -712
rect -1990 -730 -1986 -725
rect -1995 -779 -1990 -774
rect -1982 -783 -1978 -770
rect -1960 -783 -1955 -717
rect -1930 -721 -1926 -708
rect -1878 -712 -1874 -708
rect -1826 -712 -1822 -708
rect -1781 -712 -1777 -700
rect -1749 -712 -1745 -700
rect -1938 -725 -1926 -721
rect -1908 -717 -1886 -712
rect -1878 -717 -1834 -712
rect -1826 -717 -1789 -712
rect -1781 -717 -1757 -712
rect -1749 -717 -1735 -712
rect -1938 -730 -1934 -725
rect -1943 -779 -1938 -774
rect -1930 -783 -1926 -770
rect -1908 -783 -1903 -717
rect -1889 -740 -1886 -735
rect -1878 -744 -1874 -717
rect -1886 -775 -1882 -764
rect -1886 -779 -1874 -775
rect -2013 -788 -1990 -783
rect -1982 -788 -1938 -783
rect -1930 -788 -1886 -783
rect -1982 -791 -1978 -788
rect -1930 -791 -1926 -788
rect -1878 -791 -1874 -779
rect -1856 -783 -1851 -717
rect -1837 -740 -1834 -735
rect -1826 -744 -1822 -717
rect -1781 -720 -1777 -717
rect -1749 -720 -1745 -717
rect -1789 -747 -1785 -740
rect -1757 -747 -1753 -740
rect -1799 -749 -1735 -747
rect -1799 -753 -1797 -749
rect -1793 -753 -1773 -749
rect -1769 -753 -1765 -749
rect -1761 -753 -1741 -749
rect -1737 -753 -1735 -749
rect -1799 -755 -1735 -753
rect -1834 -775 -1830 -764
rect -1834 -779 -1822 -775
rect -1856 -788 -1834 -783
rect -1826 -791 -1822 -779
rect -1990 -819 -1986 -811
rect -1938 -819 -1934 -811
rect -1886 -819 -1882 -811
rect -1834 -819 -1830 -811
rect -2000 -820 -1812 -819
rect -2000 -824 -1973 -820
rect -1969 -824 -1921 -820
rect -1917 -824 -1869 -820
rect -1865 -824 -1817 -820
rect -1813 -824 -1812 -820
rect -2000 -825 -1812 -824
rect -2007 -838 -2000 -833
rect -1995 -838 -1948 -833
rect -1943 -838 -1894 -833
rect -1889 -838 -1842 -833
rect -8122 -2971 -8058 -2968
rect -8122 -2975 -8119 -2971
rect -8115 -2975 -8097 -2971
rect -8093 -2975 -8087 -2971
rect -8083 -2975 -8065 -2971
rect -8061 -2975 -8058 -2971
rect -8323 -2979 -8135 -2976
rect -8122 -2977 -8058 -2975
rect -8323 -2983 -8320 -2979
rect -8316 -2983 -8298 -2979
rect -8294 -2983 -8268 -2979
rect -8264 -2983 -8246 -2979
rect -8242 -2983 -8216 -2979
rect -8212 -2983 -8194 -2979
rect -8190 -2983 -8164 -2979
rect -8160 -2983 -8142 -2979
rect -8138 -2983 -8135 -2979
rect -8323 -2985 -8135 -2983
rect -8112 -2983 -8108 -2977
rect -8080 -2983 -8076 -2977
rect -8313 -2991 -8309 -2985
rect -8261 -2991 -8257 -2985
rect -8209 -2991 -8205 -2985
rect -8157 -2991 -8153 -2985
rect -8336 -3040 -8313 -3035
rect -8336 -3106 -8331 -3040
rect -8305 -3044 -8301 -3031
rect -8313 -3048 -8301 -3044
rect -8283 -3040 -8261 -3035
rect -8313 -3053 -8309 -3048
rect -8318 -3102 -8313 -3097
rect -8305 -3106 -8301 -3093
rect -8283 -3106 -8278 -3040
rect -8253 -3044 -8249 -3031
rect -8201 -3035 -8197 -3031
rect -8149 -3035 -8145 -3031
rect -8104 -3035 -8100 -3023
rect -8072 -3035 -8068 -3023
rect -7685 -3030 -7668 -3025
rect -7659 -3030 -6738 -3025
rect -8261 -3048 -8249 -3044
rect -8231 -3040 -8209 -3035
rect -8201 -3040 -8157 -3035
rect -8149 -3040 -8112 -3035
rect -8104 -3040 -8080 -3035
rect -8072 -3040 -7998 -3035
rect -8261 -3053 -8257 -3048
rect -8266 -3102 -8261 -3097
rect -8253 -3106 -8249 -3093
rect -8231 -3106 -8226 -3040
rect -8212 -3063 -8209 -3058
rect -8201 -3067 -8197 -3040
rect -8209 -3098 -8205 -3087
rect -8209 -3102 -8197 -3098
rect -8336 -3111 -8313 -3106
rect -8305 -3111 -8261 -3106
rect -8253 -3111 -8209 -3106
rect -8305 -3114 -8301 -3111
rect -8253 -3114 -8249 -3111
rect -8201 -3114 -8197 -3102
rect -8179 -3106 -8174 -3040
rect -8160 -3063 -8157 -3058
rect -8149 -3067 -8145 -3040
rect -8104 -3043 -8100 -3040
rect -8072 -3043 -8068 -3040
rect -8112 -3070 -8108 -3063
rect -8080 -3070 -8076 -3063
rect -8122 -3072 -8058 -3070
rect -8122 -3076 -8120 -3072
rect -8116 -3076 -8096 -3072
rect -8092 -3076 -8088 -3072
rect -8084 -3076 -8064 -3072
rect -8060 -3076 -8058 -3072
rect -8122 -3078 -8058 -3076
rect -8003 -3074 -7998 -3040
rect -7742 -3051 -7715 -3048
rect -7960 -3058 -7847 -3053
rect -7742 -3055 -7739 -3051
rect -7735 -3055 -7722 -3051
rect -7718 -3055 -7715 -3051
rect -7742 -3057 -7715 -3055
rect -7960 -3074 -7955 -3058
rect -8003 -3079 -7955 -3074
rect -8157 -3098 -8153 -3087
rect -8157 -3102 -8145 -3098
rect -8179 -3111 -8157 -3106
rect -8149 -3114 -8145 -3102
rect -8313 -3142 -8309 -3134
rect -8261 -3142 -8257 -3134
rect -8209 -3142 -8205 -3134
rect -8157 -3142 -8153 -3134
rect -8323 -3143 -8135 -3142
rect -8323 -3147 -8296 -3143
rect -8292 -3147 -8244 -3143
rect -8240 -3147 -8192 -3143
rect -8188 -3147 -8140 -3143
rect -8136 -3147 -8135 -3143
rect -8323 -3148 -8135 -3147
rect -8330 -3161 -8323 -3156
rect -8318 -3161 -8271 -3156
rect -8266 -3161 -8217 -3156
rect -8212 -3161 -8165 -3156
rect -8108 -3275 -8044 -3272
rect -8108 -3279 -8105 -3275
rect -8101 -3279 -8083 -3275
rect -8079 -3279 -8073 -3275
rect -8069 -3279 -8051 -3275
rect -8047 -3279 -8044 -3275
rect -8309 -3283 -8121 -3280
rect -8108 -3281 -8044 -3279
rect -8309 -3287 -8306 -3283
rect -8302 -3287 -8284 -3283
rect -8280 -3287 -8254 -3283
rect -8250 -3287 -8232 -3283
rect -8228 -3287 -8202 -3283
rect -8198 -3287 -8180 -3283
rect -8176 -3287 -8150 -3283
rect -8146 -3287 -8128 -3283
rect -8124 -3287 -8121 -3283
rect -8309 -3289 -8121 -3287
rect -8098 -3287 -8094 -3281
rect -8066 -3287 -8062 -3281
rect -8299 -3295 -8295 -3289
rect -8247 -3295 -8243 -3289
rect -8195 -3295 -8191 -3289
rect -8143 -3295 -8139 -3289
rect -8322 -3344 -8299 -3339
rect -8322 -3410 -8317 -3344
rect -8291 -3348 -8287 -3335
rect -8299 -3352 -8287 -3348
rect -8269 -3344 -8247 -3339
rect -8299 -3357 -8295 -3352
rect -8304 -3406 -8299 -3401
rect -8291 -3410 -8287 -3397
rect -8269 -3410 -8264 -3344
rect -8239 -3348 -8235 -3335
rect -8187 -3339 -8183 -3335
rect -8135 -3339 -8131 -3335
rect -8090 -3339 -8086 -3327
rect -8058 -3339 -8054 -3327
rect -7960 -3331 -7955 -3079
rect -7882 -3062 -7876 -3061
rect -7882 -3066 -7881 -3062
rect -7877 -3066 -7876 -3062
rect -7882 -3069 -7876 -3066
rect -7847 -3069 -7842 -3058
rect -7797 -3064 -7788 -3061
rect -7797 -3068 -7795 -3064
rect -7791 -3068 -7788 -3064
rect -7797 -3069 -7788 -3068
rect -7882 -3073 -7870 -3069
rect -7882 -3083 -7876 -3073
rect -7812 -3073 -7788 -3069
rect -7734 -3065 -7730 -3057
rect -7847 -3081 -7832 -3077
rect -7797 -3081 -7788 -3073
rect -7762 -3077 -7749 -3073
rect -7762 -3080 -7758 -3077
rect -7882 -3087 -7881 -3083
rect -7877 -3087 -7876 -3083
rect -7882 -3088 -7876 -3087
rect -7847 -3091 -7842 -3081
rect -7797 -3085 -7795 -3081
rect -7791 -3085 -7788 -3081
rect -7797 -3088 -7788 -3085
rect -7770 -3091 -7766 -3088
rect -7818 -3095 -7766 -3091
rect -7818 -3100 -7814 -3095
rect -7873 -3105 -7814 -3100
rect -7882 -3113 -7876 -3112
rect -7882 -3117 -7881 -3113
rect -7877 -3117 -7876 -3113
rect -7882 -3120 -7876 -3117
rect -7847 -3120 -7842 -3105
rect -7762 -3111 -7758 -3088
rect -7755 -3095 -7749 -3077
rect -7726 -3095 -7722 -3085
rect -7685 -3095 -7680 -3030
rect -7638 -3076 -7584 -3073
rect -7638 -3080 -7635 -3076
rect -7631 -3080 -7618 -3076
rect -7614 -3080 -7608 -3076
rect -7604 -3080 -7591 -3076
rect -7587 -3080 -7584 -3076
rect -7638 -3082 -7584 -3080
rect -7755 -3100 -7734 -3095
rect -7726 -3100 -7680 -3095
rect -7726 -3103 -7722 -3100
rect -7797 -3115 -7788 -3112
rect -7797 -3119 -7795 -3115
rect -7791 -3119 -7788 -3115
rect -7797 -3120 -7788 -3119
rect -7882 -3124 -7870 -3120
rect -7882 -3134 -7876 -3124
rect -7812 -3124 -7788 -3120
rect -7847 -3132 -7832 -3128
rect -7797 -3132 -7788 -3124
rect -7882 -3138 -7881 -3134
rect -7877 -3138 -7876 -3134
rect -7882 -3139 -7876 -3138
rect -7847 -3143 -7842 -3132
rect -7797 -3136 -7795 -3132
rect -7791 -3136 -7788 -3132
rect -7797 -3139 -7788 -3136
rect -7630 -3107 -7626 -3082
rect -7595 -3107 -7591 -3082
rect -7770 -3143 -7766 -3121
rect -7734 -3123 -7730 -3113
rect -7742 -3124 -7715 -3123
rect -7742 -3128 -7741 -3124
rect -7737 -3128 -7720 -3124
rect -7716 -3128 -7715 -3124
rect -7742 -3129 -7715 -3128
rect -7847 -3146 -7766 -3143
rect -7643 -3149 -7630 -3144
rect -7622 -3147 -7618 -3127
rect -7603 -3147 -7599 -3127
rect -7591 -3143 -7584 -3139
rect -7643 -3154 -7638 -3149
rect -7622 -3151 -7599 -3147
rect -7589 -3151 -7584 -3143
rect -7576 -3146 -7549 -3143
rect -7576 -3150 -7573 -3146
rect -7569 -3150 -7556 -3146
rect -7552 -3150 -7549 -3146
rect -7643 -3159 -7612 -3154
rect -7643 -3170 -7638 -3159
rect -7704 -3175 -7638 -3170
rect -7603 -3171 -7599 -3151
rect -7576 -3152 -7549 -3150
rect -7568 -3157 -7564 -3152
rect -7856 -3237 -7802 -3234
rect -7856 -3241 -7853 -3237
rect -7849 -3241 -7836 -3237
rect -7832 -3241 -7826 -3237
rect -7822 -3241 -7809 -3237
rect -7805 -3241 -7802 -3237
rect -7856 -3243 -7802 -3241
rect -7848 -3268 -7844 -3243
rect -7813 -3268 -7809 -3243
rect -7861 -3310 -7848 -3305
rect -7840 -3308 -7836 -3288
rect -7821 -3308 -7817 -3288
rect -7809 -3304 -7802 -3300
rect -7861 -3315 -7856 -3310
rect -7840 -3312 -7817 -3308
rect -7807 -3312 -7802 -3304
rect -7794 -3307 -7767 -3304
rect -7794 -3311 -7791 -3307
rect -7787 -3311 -7774 -3307
rect -7770 -3311 -7767 -3307
rect -7861 -3320 -7830 -3315
rect -7861 -3331 -7856 -3320
rect -7960 -3336 -7856 -3331
rect -7821 -3332 -7817 -3312
rect -7794 -3313 -7767 -3311
rect -7786 -3318 -7782 -3313
rect -7821 -3338 -7798 -3332
rect -8247 -3352 -8235 -3348
rect -8217 -3344 -8195 -3339
rect -8187 -3344 -8143 -3339
rect -8135 -3344 -8098 -3339
rect -8090 -3344 -8066 -3339
rect -8058 -3344 -8029 -3339
rect -7821 -3342 -7817 -3338
rect -8247 -3357 -8243 -3352
rect -8252 -3406 -8247 -3401
rect -8239 -3410 -8235 -3397
rect -8217 -3410 -8212 -3344
rect -8198 -3367 -8195 -3362
rect -8187 -3371 -8183 -3344
rect -8195 -3402 -8191 -3391
rect -8195 -3406 -8183 -3402
rect -8322 -3415 -8299 -3410
rect -8291 -3415 -8247 -3410
rect -8239 -3415 -8195 -3410
rect -8291 -3418 -8287 -3415
rect -8239 -3418 -8235 -3415
rect -8187 -3418 -8183 -3406
rect -8165 -3410 -8160 -3344
rect -8146 -3367 -8143 -3362
rect -8135 -3371 -8131 -3344
rect -8090 -3347 -8086 -3344
rect -8058 -3347 -8054 -3344
rect -8098 -3374 -8094 -3367
rect -8066 -3374 -8062 -3367
rect -7829 -3368 -7825 -3362
rect -7804 -3368 -7798 -3338
rect -7778 -3368 -7774 -3358
rect -7829 -3372 -7817 -3368
rect -8108 -3376 -8044 -3374
rect -8108 -3380 -8106 -3376
rect -8102 -3380 -8082 -3376
rect -8078 -3380 -8074 -3376
rect -8070 -3380 -8050 -3376
rect -8046 -3380 -8044 -3376
rect -8108 -3382 -8044 -3380
rect -7856 -3389 -7850 -3378
rect -8143 -3402 -8139 -3391
rect -7856 -3394 -7843 -3389
rect -7837 -3394 -7831 -3389
rect -7821 -3397 -7817 -3372
rect -7804 -3373 -7786 -3368
rect -7778 -3373 -7771 -3368
rect -7778 -3385 -7774 -3373
rect -8143 -3406 -8131 -3402
rect -8165 -3415 -8143 -3410
rect -8135 -3418 -8131 -3406
rect -7786 -3402 -7782 -3396
rect -7794 -3403 -7767 -3402
rect -7794 -3407 -7793 -3403
rect -7789 -3407 -7772 -3403
rect -7768 -3407 -7767 -3403
rect -7794 -3408 -7767 -3407
rect -7829 -3423 -7825 -3417
rect -7837 -3424 -7810 -3423
rect -7837 -3428 -7836 -3424
rect -7832 -3428 -7815 -3424
rect -7811 -3428 -7810 -3424
rect -7837 -3429 -7810 -3428
rect -8299 -3446 -8295 -3438
rect -8247 -3446 -8243 -3438
rect -8195 -3446 -8191 -3438
rect -8143 -3446 -8139 -3438
rect -8309 -3447 -8121 -3446
rect -8309 -3451 -8282 -3447
rect -8278 -3451 -8230 -3447
rect -8226 -3451 -8178 -3447
rect -8174 -3451 -8126 -3447
rect -8122 -3451 -8121 -3447
rect -8309 -3452 -8121 -3451
rect -8316 -3465 -8309 -3460
rect -8304 -3465 -8257 -3460
rect -8252 -3465 -8203 -3460
rect -8198 -3465 -8151 -3460
rect -7704 -3839 -7699 -3175
rect -7603 -3177 -7580 -3171
rect -7603 -3181 -7599 -3177
rect -7611 -3207 -7607 -3201
rect -7586 -3207 -7580 -3177
rect -7560 -3207 -7556 -3197
rect -7611 -3211 -7599 -3207
rect -7672 -3228 -7632 -3227
rect -7672 -3231 -7625 -3228
rect -7672 -3789 -7668 -3231
rect -7638 -3233 -7625 -3231
rect -7619 -3233 -7613 -3228
rect -7603 -3236 -7599 -3211
rect -7586 -3212 -7568 -3207
rect -7560 -3212 -7530 -3207
rect -7560 -3224 -7556 -3212
rect -7568 -3241 -7564 -3235
rect -7576 -3242 -7549 -3241
rect -7576 -3246 -7575 -3242
rect -7571 -3246 -7554 -3242
rect -7550 -3246 -7549 -3242
rect -7576 -3247 -7549 -3246
rect -7611 -3262 -7607 -3256
rect -7619 -3263 -7592 -3262
rect -7619 -3267 -7618 -3263
rect -7614 -3267 -7597 -3263
rect -7593 -3267 -7592 -3263
rect -7619 -3268 -7592 -3267
rect -7535 -3265 -7530 -3212
rect -7517 -3209 -7512 -3030
rect -7493 -3114 -7439 -3111
rect -7493 -3118 -7490 -3114
rect -7486 -3118 -7473 -3114
rect -7469 -3118 -7463 -3114
rect -7459 -3118 -7446 -3114
rect -7442 -3118 -7439 -3114
rect -7493 -3120 -7439 -3118
rect -7485 -3145 -7481 -3120
rect -7450 -3145 -7446 -3120
rect -7300 -3130 -7246 -3127
rect -7300 -3134 -7297 -3130
rect -7293 -3134 -7280 -3130
rect -7276 -3134 -7270 -3130
rect -7266 -3134 -7253 -3130
rect -7249 -3134 -7246 -3130
rect -7300 -3136 -7246 -3134
rect -7498 -3187 -7485 -3182
rect -7477 -3185 -7473 -3165
rect -7292 -3161 -7288 -3136
rect -7257 -3161 -7253 -3136
rect -7458 -3185 -7454 -3165
rect -7446 -3181 -7439 -3177
rect -7498 -3192 -7493 -3187
rect -7477 -3189 -7454 -3185
rect -7444 -3189 -7439 -3181
rect -7431 -3184 -7404 -3181
rect -7431 -3188 -7428 -3184
rect -7424 -3188 -7411 -3184
rect -7407 -3188 -7404 -3184
rect -7498 -3197 -7467 -3192
rect -7498 -3209 -7493 -3197
rect -7517 -3214 -7493 -3209
rect -7458 -3209 -7454 -3189
rect -7431 -3190 -7404 -3188
rect -7423 -3195 -7419 -3190
rect -7458 -3215 -7435 -3209
rect -7458 -3219 -7454 -3215
rect -7466 -3245 -7462 -3239
rect -7441 -3245 -7435 -3215
rect -7305 -3203 -7292 -3198
rect -7284 -3201 -7280 -3181
rect -7265 -3201 -7261 -3181
rect -7253 -3197 -7246 -3193
rect -7305 -3208 -7300 -3203
rect -7284 -3205 -7261 -3201
rect -7251 -3205 -7246 -3197
rect -7238 -3200 -7211 -3197
rect -7238 -3204 -7235 -3200
rect -7231 -3204 -7218 -3200
rect -7214 -3204 -7211 -3200
rect -7305 -3213 -7274 -3208
rect -7305 -3225 -7300 -3213
rect -7415 -3245 -7411 -3235
rect -7380 -3230 -7300 -3225
rect -7265 -3225 -7261 -3205
rect -7238 -3206 -7211 -3204
rect -7230 -3211 -7226 -3206
rect -7466 -3249 -7454 -3245
rect -7535 -3266 -7485 -3265
rect -7535 -3271 -7480 -3266
rect -7474 -3271 -7468 -3266
rect -7535 -3273 -7485 -3271
rect -7458 -3274 -7454 -3249
rect -7441 -3250 -7423 -3245
rect -7415 -3250 -7408 -3245
rect -7415 -3262 -7411 -3250
rect -7423 -3279 -7419 -3273
rect -7431 -3280 -7404 -3279
rect -7431 -3284 -7430 -3280
rect -7426 -3284 -7409 -3280
rect -7405 -3284 -7404 -3280
rect -7431 -3285 -7404 -3284
rect -7466 -3300 -7462 -3294
rect -7474 -3301 -7447 -3300
rect -7474 -3305 -7473 -3301
rect -7469 -3305 -7452 -3301
rect -7448 -3305 -7447 -3301
rect -7474 -3306 -7447 -3305
rect -7380 -3649 -7375 -3230
rect -7332 -3332 -7327 -3230
rect -7265 -3231 -7242 -3225
rect -7265 -3235 -7261 -3231
rect -7273 -3261 -7269 -3255
rect -7248 -3261 -7242 -3231
rect -7184 -3222 -7179 -3030
rect -7154 -3128 -7100 -3125
rect -7154 -3132 -7151 -3128
rect -7147 -3132 -7134 -3128
rect -7130 -3132 -7124 -3128
rect -7120 -3132 -7107 -3128
rect -7103 -3132 -7100 -3128
rect -7154 -3134 -7100 -3132
rect -7010 -3132 -6956 -3129
rect -7146 -3159 -7142 -3134
rect -7111 -3159 -7107 -3134
rect -7010 -3136 -7007 -3132
rect -7003 -3136 -6990 -3132
rect -6986 -3136 -6980 -3132
rect -6976 -3136 -6963 -3132
rect -6959 -3136 -6956 -3132
rect -7010 -3138 -6956 -3136
rect -7159 -3201 -7146 -3196
rect -7138 -3199 -7134 -3179
rect -7002 -3163 -6998 -3138
rect -6967 -3163 -6963 -3138
rect -7119 -3199 -7115 -3179
rect -7107 -3195 -7100 -3191
rect -7159 -3206 -7154 -3201
rect -7138 -3203 -7115 -3199
rect -7105 -3203 -7100 -3195
rect -7092 -3198 -7065 -3195
rect -7092 -3202 -7089 -3198
rect -7085 -3202 -7072 -3198
rect -7068 -3202 -7065 -3198
rect -7159 -3211 -7128 -3206
rect -7159 -3222 -7154 -3211
rect -7184 -3227 -7154 -3222
rect -7119 -3223 -7115 -3203
rect -7092 -3204 -7065 -3202
rect -7084 -3209 -7080 -3204
rect -7015 -3205 -7002 -3200
rect -6994 -3203 -6990 -3183
rect -6975 -3203 -6971 -3183
rect -6963 -3199 -6956 -3195
rect -7119 -3229 -7096 -3223
rect -7119 -3233 -7115 -3229
rect -7222 -3261 -7218 -3251
rect -7127 -3259 -7123 -3253
rect -7102 -3259 -7096 -3229
rect -7015 -3210 -7010 -3205
rect -6994 -3207 -6971 -3203
rect -6961 -3207 -6956 -3199
rect -6948 -3202 -6921 -3199
rect -6948 -3206 -6945 -3202
rect -6941 -3206 -6928 -3202
rect -6924 -3206 -6921 -3202
rect -7015 -3215 -6984 -3210
rect -7015 -3233 -7010 -3215
rect -6975 -3227 -6971 -3207
rect -6948 -3208 -6921 -3206
rect -6940 -3213 -6936 -3208
rect -6975 -3233 -6952 -3227
rect -6975 -3237 -6971 -3233
rect -7076 -3259 -7072 -3249
rect -7273 -3265 -7261 -3261
rect -7292 -3287 -7287 -3282
rect -7281 -3287 -7275 -3282
rect -7265 -3290 -7261 -3265
rect -7248 -3266 -7230 -3261
rect -7222 -3266 -7148 -3261
rect -7127 -3263 -7115 -3259
rect -7222 -3278 -7218 -3266
rect -7153 -3280 -7148 -3266
rect -7153 -3285 -7141 -3280
rect -7135 -3285 -7129 -3280
rect -7119 -3288 -7115 -3263
rect -7102 -3264 -7084 -3259
rect -7076 -3264 -7024 -3259
rect -7076 -3276 -7072 -3264
rect -7230 -3295 -7226 -3289
rect -7238 -3296 -7211 -3295
rect -7238 -3300 -7237 -3296
rect -7233 -3300 -7216 -3296
rect -7212 -3300 -7211 -3296
rect -7238 -3301 -7211 -3300
rect -7084 -3293 -7080 -3287
rect -7092 -3294 -7065 -3293
rect -7092 -3298 -7091 -3294
rect -7087 -3298 -7070 -3294
rect -7066 -3298 -7065 -3294
rect -7092 -3299 -7065 -3298
rect -7273 -3316 -7269 -3310
rect -7127 -3314 -7123 -3308
rect -7135 -3315 -7108 -3314
rect -7281 -3317 -7254 -3316
rect -7281 -3321 -7280 -3317
rect -7276 -3321 -7259 -3317
rect -7255 -3321 -7254 -3317
rect -7135 -3319 -7134 -3315
rect -7130 -3319 -7113 -3315
rect -7109 -3319 -7108 -3315
rect -7135 -3320 -7108 -3319
rect -7029 -3315 -7024 -3264
rect -6983 -3263 -6979 -3257
rect -6958 -3263 -6952 -3233
rect -6898 -3229 -6893 -3030
rect -6855 -3134 -6801 -3131
rect -6855 -3138 -6852 -3134
rect -6848 -3138 -6835 -3134
rect -6831 -3138 -6825 -3134
rect -6821 -3138 -6808 -3134
rect -6804 -3138 -6801 -3134
rect -6855 -3140 -6801 -3138
rect -6847 -3165 -6843 -3140
rect -6812 -3165 -6808 -3140
rect -6860 -3207 -6847 -3202
rect -6839 -3205 -6835 -3185
rect -6820 -3205 -6816 -3185
rect -6808 -3201 -6801 -3197
rect -6860 -3212 -6855 -3207
rect -6839 -3209 -6816 -3205
rect -6806 -3209 -6801 -3201
rect -6793 -3204 -6766 -3201
rect -6793 -3208 -6790 -3204
rect -6786 -3208 -6773 -3204
rect -6769 -3208 -6766 -3204
rect -6860 -3217 -6829 -3212
rect -6860 -3229 -6855 -3217
rect -6898 -3234 -6855 -3229
rect -6820 -3229 -6816 -3209
rect -6793 -3210 -6766 -3208
rect -6785 -3215 -6781 -3210
rect -6820 -3235 -6797 -3229
rect -6820 -3239 -6816 -3235
rect -6932 -3263 -6928 -3253
rect -6983 -3267 -6971 -3263
rect -7011 -3284 -7004 -3283
rect -7011 -3289 -6997 -3284
rect -6991 -3289 -6985 -3284
rect -7281 -3322 -7254 -3321
rect -7011 -3332 -7006 -3289
rect -6975 -3292 -6971 -3267
rect -6958 -3268 -6940 -3263
rect -6932 -3268 -6886 -3263
rect -6932 -3280 -6928 -3268
rect -6891 -3285 -6886 -3268
rect -6828 -3265 -6824 -3259
rect -6803 -3265 -6797 -3235
rect -6743 -3236 -6738 -3030
rect -6720 -3142 -6666 -3139
rect -6720 -3146 -6717 -3142
rect -6713 -3146 -6700 -3142
rect -6696 -3146 -6690 -3142
rect -6686 -3146 -6673 -3142
rect -6669 -3146 -6666 -3142
rect -6720 -3148 -6666 -3146
rect -6712 -3173 -6708 -3148
rect -6677 -3173 -6673 -3148
rect -6725 -3215 -6712 -3210
rect -6704 -3213 -6700 -3193
rect -6587 -3171 -6267 -3166
rect -6685 -3213 -6681 -3193
rect -6673 -3209 -6666 -3205
rect -6725 -3220 -6720 -3215
rect -6704 -3217 -6681 -3213
rect -6671 -3217 -6666 -3209
rect -6658 -3212 -6631 -3209
rect -6658 -3216 -6655 -3212
rect -6651 -3216 -6638 -3212
rect -6634 -3216 -6631 -3212
rect -6725 -3225 -6694 -3220
rect -6725 -3236 -6720 -3225
rect -6743 -3241 -6719 -3236
rect -6685 -3237 -6681 -3217
rect -6658 -3218 -6631 -3216
rect -6650 -3223 -6646 -3218
rect -6685 -3243 -6662 -3237
rect -6685 -3247 -6681 -3243
rect -6777 -3265 -6773 -3255
rect -6828 -3269 -6816 -3265
rect -6891 -3286 -6843 -3285
rect -6891 -3290 -6842 -3286
rect -6855 -3291 -6842 -3290
rect -6836 -3291 -6830 -3286
rect -6940 -3297 -6936 -3291
rect -6820 -3294 -6816 -3269
rect -6803 -3270 -6785 -3265
rect -6777 -3270 -6739 -3265
rect -6777 -3282 -6773 -3270
rect -6948 -3298 -6921 -3297
rect -6948 -3302 -6947 -3298
rect -6943 -3302 -6926 -3298
rect -6922 -3302 -6921 -3298
rect -6948 -3303 -6921 -3302
rect -6983 -3318 -6979 -3312
rect -6785 -3299 -6781 -3293
rect -6793 -3300 -6766 -3299
rect -6793 -3304 -6792 -3300
rect -6788 -3304 -6771 -3300
rect -6767 -3304 -6766 -3300
rect -6793 -3305 -6766 -3304
rect -6991 -3319 -6964 -3318
rect -6991 -3323 -6990 -3319
rect -6986 -3323 -6969 -3319
rect -6965 -3323 -6964 -3319
rect -6828 -3320 -6824 -3314
rect -6991 -3324 -6964 -3323
rect -6836 -3321 -6809 -3320
rect -6836 -3325 -6835 -3321
rect -6831 -3325 -6814 -3321
rect -6810 -3325 -6809 -3321
rect -6836 -3326 -6809 -3325
rect -7332 -3337 -7006 -3332
rect -6744 -3369 -6739 -3270
rect -6693 -3273 -6689 -3267
rect -6668 -3273 -6662 -3243
rect -6642 -3273 -6638 -3263
rect -6587 -3273 -6582 -3171
rect -6559 -3198 -6532 -3195
rect -6559 -3202 -6556 -3198
rect -6552 -3202 -6539 -3198
rect -6535 -3202 -6532 -3198
rect -6559 -3204 -6532 -3202
rect -6551 -3216 -6547 -3204
rect -6562 -3244 -6551 -3239
rect -6543 -3248 -6539 -3236
rect -6693 -3277 -6681 -3273
rect -6720 -3294 -6714 -3293
rect -6714 -3299 -6707 -3294
rect -6701 -3299 -6695 -3294
rect -6685 -3302 -6681 -3277
rect -6668 -3278 -6650 -3273
rect -6642 -3278 -6582 -3273
rect -6551 -3252 -6539 -3248
rect -6510 -3246 -6483 -3243
rect -6510 -3250 -6507 -3246
rect -6503 -3250 -6490 -3246
rect -6486 -3250 -6483 -3246
rect -6510 -3252 -6483 -3250
rect -6551 -3264 -6547 -3252
rect -6502 -3260 -6498 -3252
rect -6397 -3254 -6370 -3251
rect -6397 -3258 -6394 -3254
rect -6390 -3258 -6377 -3254
rect -6373 -3258 -6370 -3254
rect -6397 -3260 -6370 -3258
rect -6642 -3290 -6638 -3278
rect -6575 -3290 -6566 -3289
rect -6568 -3294 -6566 -3290
rect -6543 -3290 -6539 -3283
rect -6494 -3290 -6490 -3280
rect -6389 -3272 -6385 -3260
rect -6543 -3295 -6502 -3290
rect -6494 -3295 -6401 -3290
rect -6543 -3298 -6539 -3295
rect -6494 -3298 -6490 -3295
rect -6650 -3307 -6646 -3301
rect -6558 -3302 -6521 -3298
rect -6658 -3308 -6631 -3307
rect -6558 -3308 -6554 -3302
rect -6525 -3308 -6521 -3302
rect -6658 -3312 -6657 -3308
rect -6653 -3312 -6636 -3308
rect -6632 -3312 -6631 -3308
rect -6658 -3313 -6631 -3312
rect -6406 -3300 -6389 -3295
rect -6381 -3304 -6377 -3292
rect -6389 -3308 -6377 -3304
rect -6348 -3302 -6321 -3299
rect -6348 -3306 -6345 -3302
rect -6341 -3306 -6328 -3302
rect -6324 -3306 -6321 -3302
rect -6348 -3308 -6321 -3306
rect -6502 -3318 -6498 -3308
rect -6693 -3328 -6689 -3322
rect -6566 -3325 -6562 -3318
rect -6533 -3325 -6529 -3318
rect -6510 -3319 -6483 -3318
rect -6510 -3323 -6509 -3319
rect -6505 -3323 -6488 -3319
rect -6484 -3323 -6483 -3319
rect -6510 -3324 -6483 -3323
rect -6389 -3320 -6385 -3308
rect -6340 -3316 -6336 -3308
rect -6574 -3326 -6547 -3325
rect -6701 -3329 -6674 -3328
rect -6701 -3333 -6700 -3329
rect -6696 -3333 -6679 -3329
rect -6675 -3333 -6674 -3329
rect -6574 -3330 -6573 -3326
rect -6569 -3330 -6552 -3326
rect -6548 -3330 -6547 -3326
rect -6574 -3331 -6547 -3330
rect -6541 -3326 -6514 -3325
rect -6541 -3330 -6540 -3326
rect -6536 -3330 -6519 -3326
rect -6515 -3330 -6514 -3326
rect -6541 -3331 -6514 -3330
rect -6701 -3334 -6674 -3333
rect -6272 -3328 -6267 -3171
rect -6239 -3310 -6212 -3307
rect -6239 -3314 -6236 -3310
rect -6232 -3314 -6219 -3310
rect -6215 -3314 -6212 -3310
rect -6239 -3316 -6212 -3314
rect -6231 -3328 -6227 -3316
rect -6429 -3350 -6404 -3345
rect -6381 -3346 -6377 -3339
rect -6332 -3346 -6328 -3336
rect -6429 -3369 -6424 -3350
rect -6381 -3351 -6340 -3346
rect -6332 -3351 -6251 -3346
rect -6381 -3354 -6377 -3351
rect -6332 -3354 -6328 -3351
rect -6396 -3358 -6359 -3354
rect -6396 -3364 -6392 -3358
rect -6363 -3364 -6359 -3358
rect -6744 -3374 -6424 -3369
rect -6256 -3356 -6231 -3351
rect -6223 -3360 -6219 -3348
rect -6231 -3364 -6219 -3360
rect -6190 -3358 -6163 -3355
rect -6190 -3362 -6187 -3358
rect -6183 -3362 -6170 -3358
rect -6166 -3362 -6163 -3358
rect -6190 -3364 -6163 -3362
rect -6340 -3374 -6336 -3364
rect -6404 -3381 -6400 -3374
rect -6371 -3381 -6367 -3374
rect -6348 -3375 -6321 -3374
rect -6348 -3379 -6347 -3375
rect -6343 -3379 -6326 -3375
rect -6322 -3379 -6321 -3375
rect -6348 -3380 -6321 -3379
rect -6231 -3376 -6227 -3364
rect -6182 -3372 -6178 -3364
rect -6412 -3382 -6385 -3381
rect -6412 -3386 -6411 -3382
rect -6407 -3386 -6390 -3382
rect -6386 -3386 -6385 -3382
rect -6412 -3387 -6385 -3386
rect -6379 -3382 -6352 -3381
rect -6379 -3386 -6378 -3382
rect -6374 -3386 -6357 -3382
rect -6353 -3386 -6352 -3382
rect -6379 -3387 -6352 -3386
rect -6073 -3386 -6046 -3383
rect -6073 -3390 -6070 -3386
rect -6066 -3390 -6053 -3386
rect -6049 -3390 -6046 -3386
rect -6073 -3392 -6046 -3390
rect -6251 -3405 -6246 -3401
rect -6255 -3406 -6246 -3405
rect -6223 -3402 -6219 -3395
rect -6174 -3402 -6170 -3392
rect -6223 -3407 -6182 -3402
rect -6174 -3407 -6083 -3402
rect -6223 -3410 -6219 -3407
rect -6174 -3410 -6170 -3407
rect -6238 -3414 -6201 -3410
rect -6238 -3420 -6234 -3414
rect -6205 -3420 -6201 -3414
rect -6182 -3430 -6178 -3420
rect -6088 -3427 -6083 -3407
rect -6065 -3404 -6061 -3392
rect -6246 -3437 -6242 -3430
rect -6213 -3437 -6209 -3430
rect -6190 -3431 -6163 -3430
rect -6190 -3435 -6189 -3431
rect -6185 -3435 -6168 -3431
rect -6164 -3435 -6163 -3431
rect -6088 -3432 -6065 -3427
rect -6190 -3436 -6163 -3435
rect -6057 -3436 -6053 -3424
rect -5722 -3425 -5658 -3422
rect -5722 -3429 -5719 -3425
rect -5715 -3429 -5697 -3425
rect -5693 -3429 -5687 -3425
rect -5683 -3429 -5665 -3425
rect -5661 -3429 -5658 -3425
rect -6254 -3438 -6227 -3437
rect -6254 -3442 -6253 -3438
rect -6249 -3442 -6232 -3438
rect -6228 -3442 -6227 -3438
rect -6254 -3443 -6227 -3442
rect -6221 -3438 -6194 -3437
rect -6221 -3442 -6220 -3438
rect -6216 -3442 -6199 -3438
rect -6195 -3442 -6194 -3438
rect -6221 -3443 -6194 -3442
rect -6065 -3440 -6053 -3436
rect -6024 -3434 -5997 -3431
rect -6024 -3438 -6021 -3434
rect -6017 -3438 -6004 -3434
rect -6000 -3438 -5997 -3434
rect -6024 -3440 -5997 -3438
rect -5923 -3433 -5735 -3430
rect -5722 -3431 -5658 -3429
rect -5923 -3437 -5920 -3433
rect -5916 -3437 -5898 -3433
rect -5894 -3437 -5868 -3433
rect -5864 -3437 -5846 -3433
rect -5842 -3437 -5816 -3433
rect -5812 -3437 -5794 -3433
rect -5790 -3437 -5764 -3433
rect -5760 -3437 -5742 -3433
rect -5738 -3437 -5735 -3433
rect -5923 -3439 -5735 -3437
rect -5712 -3437 -5708 -3431
rect -5680 -3437 -5676 -3431
rect -6065 -3452 -6061 -3440
rect -6016 -3448 -6012 -3440
rect -5913 -3445 -5909 -3439
rect -5861 -3445 -5857 -3439
rect -5809 -3445 -5805 -3439
rect -5757 -3445 -5753 -3439
rect -6083 -3482 -6080 -3477
rect -6057 -3478 -6053 -3471
rect -6008 -3478 -6004 -3468
rect -6057 -3483 -6016 -3478
rect -6008 -3483 -5931 -3478
rect -6057 -3486 -6053 -3483
rect -6008 -3486 -6004 -3483
rect -6072 -3490 -6035 -3486
rect -6072 -3496 -6068 -3490
rect -6039 -3496 -6035 -3490
rect -5936 -3489 -5931 -3483
rect -5553 -3467 -5526 -3464
rect -5553 -3471 -5550 -3467
rect -5546 -3471 -5533 -3467
rect -5529 -3471 -5526 -3467
rect -5553 -3473 -5526 -3471
rect -5936 -3494 -5913 -3489
rect -6016 -3506 -6012 -3496
rect -6080 -3513 -6076 -3506
rect -6047 -3513 -6043 -3506
rect -6024 -3507 -5997 -3506
rect -6024 -3511 -6023 -3507
rect -6019 -3511 -6002 -3507
rect -5998 -3511 -5997 -3507
rect -6024 -3512 -5997 -3511
rect -6088 -3514 -6061 -3513
rect -6088 -3518 -6087 -3514
rect -6083 -3518 -6066 -3514
rect -6062 -3518 -6061 -3514
rect -6088 -3519 -6061 -3518
rect -6055 -3514 -6028 -3513
rect -6055 -3518 -6054 -3514
rect -6050 -3518 -6033 -3514
rect -6029 -3518 -6028 -3514
rect -6055 -3519 -6028 -3518
rect -5936 -3560 -5931 -3494
rect -5905 -3498 -5901 -3485
rect -5913 -3502 -5901 -3498
rect -5883 -3494 -5861 -3489
rect -5913 -3507 -5909 -3502
rect -5918 -3556 -5913 -3551
rect -5905 -3560 -5901 -3547
rect -5883 -3560 -5878 -3494
rect -5853 -3498 -5849 -3485
rect -5801 -3489 -5797 -3485
rect -5749 -3489 -5745 -3485
rect -5704 -3489 -5700 -3477
rect -5672 -3489 -5668 -3477
rect -5545 -3478 -5541 -3473
rect -5861 -3502 -5849 -3498
rect -5831 -3494 -5809 -3489
rect -5801 -3494 -5757 -3489
rect -5749 -3494 -5712 -3489
rect -5704 -3494 -5680 -3489
rect -5672 -3494 -5569 -3489
rect -5861 -3507 -5857 -3502
rect -5866 -3556 -5861 -3551
rect -5853 -3560 -5849 -3547
rect -5831 -3560 -5826 -3494
rect -5812 -3517 -5809 -3512
rect -5801 -3521 -5797 -3494
rect -5809 -3552 -5805 -3541
rect -5809 -3556 -5797 -3552
rect -5936 -3565 -5913 -3560
rect -5905 -3565 -5861 -3560
rect -5853 -3565 -5809 -3560
rect -5905 -3568 -5901 -3565
rect -5853 -3568 -5849 -3565
rect -5801 -3568 -5797 -3556
rect -5779 -3560 -5774 -3494
rect -5760 -3517 -5757 -3512
rect -5749 -3521 -5745 -3494
rect -5704 -3497 -5700 -3494
rect -5672 -3497 -5668 -3494
rect -5712 -3524 -5708 -3517
rect -5680 -3524 -5676 -3517
rect -5722 -3526 -5658 -3524
rect -5722 -3530 -5720 -3526
rect -5716 -3530 -5696 -3526
rect -5692 -3530 -5688 -3526
rect -5684 -3530 -5664 -3526
rect -5660 -3530 -5658 -3526
rect -5722 -3532 -5658 -3530
rect -5574 -3528 -5569 -3494
rect -5537 -3528 -5533 -3518
rect -5574 -3533 -5545 -3528
rect -5537 -3533 -5524 -3528
rect -5757 -3552 -5753 -3541
rect -5537 -3545 -5533 -3533
rect -5757 -3556 -5745 -3552
rect -5779 -3565 -5757 -3560
rect -5749 -3568 -5745 -3556
rect -5545 -3562 -5541 -3556
rect -5553 -3563 -5526 -3562
rect -5553 -3567 -5552 -3563
rect -5548 -3567 -5531 -3563
rect -5527 -3567 -5526 -3563
rect -5553 -3568 -5526 -3567
rect -5913 -3596 -5909 -3588
rect -5861 -3596 -5857 -3588
rect -5809 -3596 -5805 -3588
rect -5757 -3596 -5753 -3588
rect -5923 -3597 -5735 -3596
rect -5923 -3601 -5896 -3597
rect -5892 -3601 -5844 -3597
rect -5840 -3601 -5792 -3597
rect -5788 -3601 -5740 -3597
rect -5736 -3601 -5735 -3597
rect -5923 -3602 -5735 -3601
rect -5930 -3615 -5923 -3610
rect -5918 -3615 -5871 -3610
rect -5866 -3615 -5817 -3610
rect -5812 -3615 -5765 -3610
rect -7380 -3654 -7079 -3649
rect -7672 -3793 -7356 -3789
rect -7704 -3844 -7670 -3839
rect -7675 -3874 -7670 -3844
rect -7360 -3862 -7356 -3793
rect -7360 -3866 -7355 -3862
rect -7084 -3874 -7079 -3654
rect -7066 -3765 -6303 -3760
rect -7675 -3879 -7026 -3874
rect -8053 -3883 -7989 -3880
rect -8053 -3887 -8050 -3883
rect -8046 -3887 -8028 -3883
rect -8024 -3887 -8018 -3883
rect -8014 -3887 -7996 -3883
rect -7992 -3887 -7989 -3883
rect -8254 -3891 -8066 -3888
rect -8053 -3889 -7989 -3887
rect -8254 -3895 -8251 -3891
rect -8247 -3895 -8229 -3891
rect -8225 -3895 -8199 -3891
rect -8195 -3895 -8177 -3891
rect -8173 -3895 -8147 -3891
rect -8143 -3895 -8125 -3891
rect -8121 -3895 -8095 -3891
rect -8091 -3895 -8073 -3891
rect -8069 -3895 -8066 -3891
rect -8254 -3897 -8066 -3895
rect -8043 -3895 -8039 -3889
rect -8011 -3895 -8007 -3889
rect -8244 -3903 -8240 -3897
rect -8192 -3903 -8188 -3897
rect -8140 -3903 -8136 -3897
rect -8088 -3903 -8084 -3897
rect -7736 -3902 -7709 -3899
rect -8267 -3952 -8244 -3947
rect -8267 -4018 -8262 -3952
rect -8236 -3956 -8232 -3943
rect -8244 -3960 -8232 -3956
rect -8214 -3952 -8192 -3947
rect -8244 -3965 -8240 -3960
rect -8249 -4014 -8244 -4009
rect -8236 -4018 -8232 -4005
rect -8214 -4018 -8209 -3952
rect -8184 -3956 -8180 -3943
rect -8132 -3947 -8128 -3943
rect -8080 -3947 -8076 -3943
rect -8035 -3947 -8031 -3935
rect -8003 -3947 -7999 -3935
rect -7904 -3909 -7841 -3904
rect -7736 -3906 -7733 -3902
rect -7729 -3906 -7716 -3902
rect -7712 -3906 -7709 -3902
rect -7736 -3908 -7709 -3906
rect -7904 -3947 -7899 -3909
rect -7876 -3913 -7870 -3912
rect -7876 -3917 -7875 -3913
rect -7871 -3917 -7870 -3913
rect -7876 -3920 -7870 -3917
rect -7841 -3920 -7836 -3909
rect -7791 -3915 -7782 -3912
rect -7791 -3919 -7789 -3915
rect -7785 -3919 -7782 -3915
rect -7791 -3920 -7782 -3919
rect -7876 -3924 -7864 -3920
rect -7876 -3934 -7870 -3924
rect -7806 -3924 -7782 -3920
rect -7728 -3916 -7724 -3908
rect -7841 -3932 -7826 -3928
rect -7791 -3932 -7782 -3924
rect -7756 -3928 -7743 -3924
rect -7756 -3931 -7752 -3928
rect -7876 -3938 -7875 -3934
rect -7871 -3938 -7870 -3934
rect -7876 -3939 -7870 -3938
rect -7841 -3942 -7836 -3932
rect -7791 -3936 -7789 -3932
rect -7785 -3936 -7782 -3932
rect -7791 -3939 -7782 -3936
rect -7764 -3942 -7760 -3939
rect -7812 -3946 -7760 -3942
rect -8192 -3960 -8180 -3956
rect -8162 -3952 -8140 -3947
rect -8132 -3952 -8088 -3947
rect -8080 -3952 -8043 -3947
rect -8035 -3952 -8011 -3947
rect -8003 -3952 -7899 -3947
rect -7812 -3951 -7808 -3946
rect -8192 -3965 -8188 -3960
rect -8197 -4014 -8192 -4009
rect -8184 -4018 -8180 -4005
rect -8162 -4018 -8157 -3952
rect -8143 -3975 -8140 -3970
rect -8132 -3979 -8128 -3952
rect -8140 -4010 -8136 -3999
rect -8140 -4014 -8128 -4010
rect -8267 -4023 -8244 -4018
rect -8236 -4023 -8192 -4018
rect -8184 -4023 -8140 -4018
rect -8236 -4026 -8232 -4023
rect -8184 -4026 -8180 -4023
rect -8132 -4026 -8128 -4014
rect -8110 -4018 -8105 -3952
rect -8091 -3975 -8088 -3970
rect -8080 -3979 -8076 -3952
rect -8035 -3955 -8031 -3952
rect -8003 -3955 -7999 -3952
rect -8043 -3982 -8039 -3975
rect -8011 -3982 -8007 -3975
rect -8053 -3984 -7989 -3982
rect -8053 -3988 -8051 -3984
rect -8047 -3988 -8027 -3984
rect -8023 -3988 -8019 -3984
rect -8015 -3988 -7995 -3984
rect -7991 -3988 -7989 -3984
rect -8053 -3990 -7989 -3988
rect -8088 -4010 -8084 -3999
rect -8088 -4014 -8076 -4010
rect -8110 -4023 -8088 -4018
rect -8080 -4026 -8076 -4014
rect -8244 -4054 -8240 -4046
rect -8192 -4054 -8188 -4046
rect -8140 -4054 -8136 -4046
rect -8088 -4054 -8084 -4046
rect -8254 -4055 -8066 -4054
rect -8254 -4059 -8227 -4055
rect -8223 -4059 -8175 -4055
rect -8171 -4059 -8123 -4055
rect -8119 -4059 -8071 -4055
rect -8067 -4059 -8066 -4055
rect -8254 -4060 -8066 -4059
rect -8261 -4073 -8254 -4068
rect -8249 -4073 -8202 -4068
rect -8197 -4073 -8148 -4068
rect -8143 -4073 -8096 -4068
rect -8036 -4124 -7972 -4121
rect -8036 -4128 -8033 -4124
rect -8029 -4128 -8011 -4124
rect -8007 -4128 -8001 -4124
rect -7997 -4128 -7979 -4124
rect -7975 -4128 -7972 -4124
rect -8237 -4132 -8049 -4129
rect -8036 -4130 -7972 -4128
rect -8237 -4136 -8234 -4132
rect -8230 -4136 -8212 -4132
rect -8208 -4136 -8182 -4132
rect -8178 -4136 -8160 -4132
rect -8156 -4136 -8130 -4132
rect -8126 -4136 -8108 -4132
rect -8104 -4136 -8078 -4132
rect -8074 -4136 -8056 -4132
rect -8052 -4136 -8049 -4132
rect -8237 -4138 -8049 -4136
rect -8026 -4136 -8022 -4130
rect -7994 -4136 -7990 -4130
rect -8227 -4144 -8223 -4138
rect -8175 -4144 -8171 -4138
rect -8123 -4144 -8119 -4138
rect -8071 -4144 -8067 -4138
rect -8250 -4193 -8227 -4188
rect -8250 -4259 -8245 -4193
rect -8219 -4197 -8215 -4184
rect -8227 -4201 -8215 -4197
rect -8197 -4193 -8175 -4188
rect -8227 -4206 -8223 -4201
rect -8232 -4255 -8227 -4250
rect -8219 -4259 -8215 -4246
rect -8197 -4259 -8192 -4193
rect -8167 -4197 -8163 -4184
rect -8115 -4188 -8111 -4184
rect -8063 -4188 -8059 -4184
rect -8018 -4188 -8014 -4176
rect -7986 -4188 -7982 -4176
rect -8175 -4201 -8163 -4197
rect -8145 -4193 -8123 -4188
rect -8115 -4193 -8071 -4188
rect -8063 -4193 -8026 -4188
rect -8018 -4193 -7994 -4188
rect -7986 -4193 -7931 -4188
rect -8175 -4206 -8171 -4201
rect -8180 -4255 -8175 -4250
rect -8167 -4259 -8163 -4246
rect -8145 -4259 -8140 -4193
rect -8126 -4216 -8123 -4211
rect -8115 -4220 -8111 -4193
rect -8123 -4251 -8119 -4240
rect -8123 -4255 -8111 -4251
rect -8250 -4264 -8227 -4259
rect -8219 -4264 -8175 -4259
rect -8167 -4264 -8123 -4259
rect -8219 -4267 -8215 -4264
rect -8167 -4267 -8163 -4264
rect -8115 -4267 -8111 -4255
rect -8093 -4259 -8088 -4193
rect -8074 -4216 -8071 -4211
rect -8063 -4220 -8059 -4193
rect -8018 -4196 -8014 -4193
rect -7986 -4196 -7982 -4193
rect -8026 -4223 -8022 -4216
rect -7994 -4223 -7990 -4216
rect -8036 -4225 -7972 -4223
rect -8036 -4229 -8034 -4225
rect -8030 -4229 -8010 -4225
rect -8006 -4229 -8002 -4225
rect -7998 -4229 -7978 -4225
rect -7974 -4229 -7972 -4225
rect -8036 -4231 -7972 -4229
rect -8071 -4251 -8067 -4240
rect -8071 -4255 -8059 -4251
rect -8093 -4264 -8071 -4259
rect -8063 -4267 -8059 -4255
rect -7936 -4274 -7931 -4193
rect -7904 -4247 -7899 -3952
rect -7871 -3956 -7808 -3951
rect -7876 -3964 -7870 -3963
rect -7876 -3968 -7875 -3964
rect -7871 -3968 -7870 -3964
rect -7876 -3971 -7870 -3968
rect -7841 -3971 -7836 -3956
rect -7756 -3962 -7752 -3939
rect -7749 -3946 -7743 -3928
rect -7720 -3946 -7716 -3936
rect -7675 -3946 -7670 -3879
rect -7630 -3891 -7576 -3888
rect -7630 -3895 -7627 -3891
rect -7623 -3895 -7610 -3891
rect -7606 -3895 -7600 -3891
rect -7596 -3895 -7583 -3891
rect -7579 -3895 -7576 -3891
rect -7630 -3897 -7576 -3895
rect -7461 -3890 -7407 -3887
rect -7461 -3894 -7458 -3890
rect -7454 -3894 -7441 -3890
rect -7437 -3894 -7431 -3890
rect -7427 -3894 -7414 -3890
rect -7410 -3894 -7407 -3890
rect -7461 -3896 -7407 -3894
rect -7622 -3922 -7618 -3897
rect -7587 -3922 -7583 -3897
rect -7749 -3951 -7728 -3946
rect -7720 -3951 -7670 -3946
rect -7720 -3954 -7716 -3951
rect -7791 -3966 -7782 -3963
rect -7791 -3970 -7789 -3966
rect -7785 -3970 -7782 -3966
rect -7791 -3971 -7782 -3970
rect -7876 -3975 -7864 -3971
rect -7876 -3985 -7870 -3975
rect -7806 -3975 -7782 -3971
rect -7841 -3983 -7826 -3979
rect -7791 -3983 -7782 -3975
rect -7876 -3989 -7875 -3985
rect -7871 -3989 -7870 -3985
rect -7876 -3990 -7870 -3989
rect -7841 -3994 -7836 -3983
rect -7791 -3987 -7789 -3983
rect -7785 -3987 -7782 -3983
rect -7791 -3990 -7782 -3987
rect -7764 -3994 -7760 -3972
rect -7728 -3974 -7724 -3964
rect -7736 -3975 -7709 -3974
rect -7736 -3979 -7735 -3975
rect -7731 -3979 -7714 -3975
rect -7710 -3979 -7709 -3975
rect -7736 -3980 -7709 -3979
rect -7841 -3997 -7760 -3994
rect -7863 -4152 -7809 -4149
rect -7863 -4156 -7860 -4152
rect -7856 -4156 -7843 -4152
rect -7839 -4156 -7833 -4152
rect -7829 -4156 -7816 -4152
rect -7812 -4156 -7809 -4152
rect -7863 -4158 -7809 -4156
rect -7855 -4183 -7851 -4158
rect -7820 -4183 -7816 -4158
rect -7868 -4225 -7855 -4220
rect -7847 -4223 -7843 -4203
rect -7828 -4223 -7824 -4203
rect -7816 -4219 -7809 -4215
rect -7868 -4230 -7863 -4225
rect -7847 -4227 -7824 -4223
rect -7814 -4227 -7809 -4219
rect -7801 -4222 -7774 -4219
rect -7801 -4226 -7798 -4222
rect -7794 -4226 -7781 -4222
rect -7777 -4226 -7774 -4222
rect -7868 -4235 -7837 -4230
rect -7868 -4247 -7863 -4235
rect -7904 -4252 -7863 -4247
rect -7828 -4247 -7824 -4227
rect -7801 -4228 -7774 -4226
rect -7793 -4233 -7789 -4228
rect -7828 -4253 -7805 -4247
rect -7828 -4257 -7824 -4253
rect -7936 -4279 -7890 -4274
rect -7836 -4283 -7832 -4277
rect -7811 -4283 -7805 -4253
rect -7675 -4254 -7670 -3951
rect -7635 -3964 -7622 -3959
rect -7614 -3962 -7610 -3942
rect -7453 -3921 -7449 -3896
rect -7418 -3921 -7414 -3896
rect -7595 -3962 -7591 -3942
rect -7583 -3958 -7576 -3954
rect -7635 -3969 -7630 -3964
rect -7614 -3966 -7591 -3962
rect -7581 -3966 -7576 -3958
rect -7568 -3961 -7541 -3958
rect -7568 -3965 -7565 -3961
rect -7561 -3965 -7548 -3961
rect -7544 -3965 -7541 -3961
rect -7635 -3974 -7604 -3969
rect -7635 -3990 -7630 -3974
rect -7595 -3986 -7591 -3966
rect -7568 -3967 -7541 -3965
rect -7466 -3963 -7453 -3958
rect -7445 -3961 -7441 -3941
rect -7426 -3961 -7422 -3941
rect -7414 -3957 -7407 -3953
rect -7560 -3972 -7556 -3967
rect -7466 -3968 -7461 -3963
rect -7445 -3965 -7422 -3961
rect -7412 -3965 -7407 -3957
rect -7399 -3960 -7372 -3957
rect -7399 -3964 -7396 -3960
rect -7392 -3964 -7379 -3960
rect -7375 -3964 -7372 -3960
rect -7595 -3992 -7572 -3986
rect -7595 -3996 -7591 -3992
rect -7603 -4022 -7599 -4016
rect -7578 -4022 -7572 -3992
rect -7466 -3973 -7435 -3968
rect -7466 -3983 -7461 -3973
rect -7426 -3985 -7422 -3965
rect -7399 -3966 -7372 -3964
rect -7391 -3971 -7387 -3966
rect -7426 -3991 -7403 -3985
rect -7426 -3995 -7422 -3991
rect -7552 -4022 -7548 -4012
rect -7434 -4021 -7430 -4015
rect -7409 -4021 -7403 -3991
rect -7383 -4021 -7379 -4011
rect -7360 -4021 -7355 -3901
rect -7334 -3981 -7329 -3879
rect -7297 -3888 -7243 -3885
rect -7297 -3892 -7294 -3888
rect -7290 -3892 -7277 -3888
rect -7273 -3892 -7267 -3888
rect -7263 -3892 -7250 -3888
rect -7246 -3892 -7243 -3888
rect -7297 -3894 -7243 -3892
rect -7157 -3890 -7103 -3887
rect -7157 -3894 -7154 -3890
rect -7150 -3894 -7137 -3890
rect -7133 -3894 -7127 -3890
rect -7123 -3894 -7110 -3890
rect -7106 -3894 -7103 -3890
rect -7289 -3919 -7285 -3894
rect -7254 -3919 -7250 -3894
rect -7157 -3896 -7103 -3894
rect -7302 -3961 -7289 -3956
rect -7281 -3959 -7277 -3939
rect -7149 -3921 -7145 -3896
rect -7114 -3921 -7110 -3896
rect -7262 -3959 -7258 -3939
rect -7250 -3955 -7243 -3951
rect -7302 -3966 -7297 -3961
rect -7281 -3963 -7258 -3959
rect -7248 -3963 -7243 -3955
rect -7235 -3958 -7208 -3955
rect -7235 -3962 -7232 -3958
rect -7228 -3962 -7215 -3958
rect -7211 -3962 -7208 -3958
rect -7302 -3971 -7271 -3966
rect -7302 -3981 -7297 -3971
rect -7334 -3986 -7297 -3981
rect -7262 -3983 -7258 -3963
rect -7235 -3964 -7208 -3962
rect -7162 -3963 -7149 -3958
rect -7141 -3961 -7137 -3941
rect -7122 -3961 -7118 -3941
rect -7110 -3957 -7103 -3953
rect -7227 -3969 -7223 -3964
rect -7162 -3968 -7157 -3963
rect -7141 -3965 -7118 -3961
rect -7108 -3965 -7103 -3957
rect -7095 -3960 -7068 -3957
rect -7095 -3964 -7092 -3960
rect -7088 -3964 -7075 -3960
rect -7071 -3964 -7068 -3960
rect -7262 -3989 -7239 -3983
rect -7262 -3993 -7258 -3989
rect -7270 -4019 -7266 -4013
rect -7245 -4019 -7239 -3989
rect -7162 -3973 -7131 -3968
rect -7162 -3984 -7157 -3973
rect -7169 -3989 -7157 -3984
rect -7122 -3985 -7118 -3965
rect -7095 -3966 -7068 -3964
rect -7087 -3971 -7083 -3966
rect -7122 -3991 -7099 -3985
rect -7122 -3995 -7118 -3991
rect -7219 -4019 -7215 -4009
rect -7603 -4026 -7591 -4022
rect -7621 -4048 -7617 -4043
rect -7611 -4048 -7605 -4043
rect -7595 -4051 -7591 -4026
rect -7578 -4027 -7560 -4022
rect -7552 -4027 -7455 -4022
rect -7434 -4025 -7422 -4021
rect -7552 -4039 -7548 -4027
rect -7461 -4042 -7455 -4027
rect -7461 -4047 -7448 -4042
rect -7442 -4047 -7436 -4042
rect -7426 -4050 -7422 -4025
rect -7409 -4026 -7391 -4021
rect -7383 -4026 -7291 -4021
rect -7270 -4023 -7258 -4019
rect -7383 -4038 -7379 -4026
rect -7560 -4056 -7556 -4050
rect -7568 -4057 -7541 -4056
rect -7568 -4061 -7567 -4057
rect -7563 -4061 -7546 -4057
rect -7542 -4061 -7541 -4057
rect -7568 -4062 -7541 -4061
rect -7297 -4040 -7291 -4026
rect -7297 -4045 -7284 -4040
rect -7278 -4045 -7272 -4040
rect -7262 -4048 -7258 -4023
rect -7245 -4024 -7227 -4019
rect -7219 -4024 -7179 -4019
rect -7219 -4036 -7215 -4024
rect -7391 -4055 -7387 -4049
rect -7399 -4056 -7372 -4055
rect -7399 -4060 -7398 -4056
rect -7394 -4060 -7377 -4056
rect -7373 -4060 -7372 -4056
rect -7399 -4061 -7372 -4060
rect -7227 -4053 -7223 -4047
rect -7235 -4054 -7208 -4053
rect -7235 -4058 -7234 -4054
rect -7230 -4058 -7213 -4054
rect -7209 -4058 -7208 -4054
rect -7235 -4059 -7208 -4058
rect -7603 -4077 -7599 -4071
rect -7434 -4076 -7430 -4070
rect -7270 -4074 -7266 -4068
rect -7278 -4075 -7251 -4074
rect -7442 -4077 -7415 -4076
rect -7611 -4078 -7584 -4077
rect -7611 -4082 -7610 -4078
rect -7606 -4082 -7589 -4078
rect -7585 -4082 -7584 -4078
rect -7442 -4081 -7441 -4077
rect -7437 -4081 -7420 -4077
rect -7416 -4081 -7415 -4077
rect -7278 -4079 -7277 -4075
rect -7273 -4079 -7256 -4075
rect -7252 -4079 -7251 -4075
rect -7278 -4080 -7251 -4079
rect -7442 -4082 -7415 -4081
rect -7611 -4083 -7584 -4082
rect -7184 -4252 -7179 -4024
rect -7130 -4021 -7126 -4015
rect -7105 -4021 -7099 -3991
rect -7031 -3997 -7026 -3879
rect -7006 -3903 -6952 -3900
rect -7006 -3907 -7003 -3903
rect -6999 -3907 -6986 -3903
rect -6982 -3907 -6976 -3903
rect -6972 -3907 -6959 -3903
rect -6955 -3907 -6952 -3903
rect -7006 -3909 -6952 -3907
rect -6998 -3934 -6994 -3909
rect -6963 -3934 -6959 -3909
rect -7011 -3976 -6998 -3971
rect -6990 -3974 -6986 -3954
rect -6696 -3945 -6669 -3942
rect -6696 -3949 -6693 -3945
rect -6689 -3949 -6676 -3945
rect -6672 -3949 -6669 -3945
rect -6696 -3951 -6669 -3949
rect -6971 -3974 -6967 -3954
rect -6688 -3963 -6684 -3951
rect -6959 -3970 -6952 -3966
rect -7011 -3981 -7006 -3976
rect -6990 -3978 -6967 -3974
rect -6957 -3978 -6952 -3970
rect -6944 -3973 -6917 -3970
rect -6944 -3977 -6941 -3973
rect -6937 -3977 -6924 -3973
rect -6920 -3977 -6917 -3973
rect -7011 -3986 -6980 -3981
rect -7011 -3997 -7006 -3986
rect -7031 -4002 -7006 -3997
rect -6971 -3998 -6967 -3978
rect -6944 -3979 -6917 -3977
rect -6936 -3984 -6932 -3979
rect -6971 -4004 -6948 -3998
rect -6971 -4008 -6967 -4004
rect -7079 -4021 -7075 -4011
rect -7130 -4025 -7118 -4021
rect -7148 -4047 -7144 -4042
rect -7138 -4047 -7132 -4042
rect -7122 -4050 -7118 -4025
rect -7105 -4026 -7087 -4021
rect -7079 -4026 -7048 -4021
rect -7041 -4026 -7000 -4021
rect -7079 -4038 -7075 -4026
rect -7087 -4055 -7083 -4049
rect -7005 -4054 -7000 -4026
rect -6979 -4034 -6975 -4028
rect -6954 -4034 -6948 -4004
rect -6928 -4034 -6924 -4024
rect -6907 -3986 -6709 -3983
rect -6907 -3988 -6688 -3986
rect -6907 -4034 -6902 -3988
rect -6979 -4038 -6967 -4034
rect -7006 -4055 -7000 -4054
rect -7095 -4056 -7068 -4055
rect -7095 -4060 -7094 -4056
rect -7090 -4060 -7073 -4056
rect -7069 -4060 -7068 -4056
rect -7006 -4060 -6993 -4055
rect -6987 -4060 -6981 -4055
rect -7095 -4061 -7068 -4060
rect -6971 -4063 -6967 -4038
rect -6954 -4039 -6936 -4034
rect -6928 -4039 -6902 -4034
rect -6928 -4051 -6924 -4039
rect -7130 -4076 -7126 -4070
rect -7138 -4077 -7111 -4076
rect -7138 -4081 -7137 -4077
rect -7133 -4081 -7116 -4077
rect -7112 -4081 -7111 -4077
rect -7138 -4082 -7111 -4081
rect -6936 -4068 -6932 -4062
rect -6944 -4069 -6917 -4068
rect -6944 -4073 -6943 -4069
rect -6939 -4073 -6922 -4069
rect -6918 -4073 -6917 -4069
rect -6944 -4074 -6917 -4073
rect -6979 -4089 -6975 -4083
rect -6987 -4090 -6960 -4089
rect -6987 -4094 -6986 -4090
rect -6982 -4094 -6965 -4090
rect -6961 -4094 -6960 -4090
rect -6987 -4095 -6960 -4094
rect -6882 -4202 -6877 -3988
rect -6714 -3991 -6688 -3988
rect -6680 -3995 -6676 -3983
rect -6688 -3999 -6676 -3995
rect -6647 -3993 -6620 -3990
rect -6647 -3997 -6644 -3993
rect -6640 -3997 -6627 -3993
rect -6623 -3997 -6620 -3993
rect -6647 -3999 -6620 -3997
rect -6688 -4011 -6684 -3999
rect -6639 -4007 -6635 -3999
rect -6708 -4041 -6703 -4036
rect -6680 -4037 -6676 -4030
rect -6631 -4037 -6627 -4027
rect -6680 -4042 -6639 -4037
rect -6631 -4042 -6608 -4037
rect -6680 -4045 -6676 -4042
rect -6631 -4045 -6627 -4042
rect -6695 -4049 -6658 -4045
rect -6695 -4055 -6691 -4049
rect -6662 -4055 -6658 -4049
rect -6639 -4065 -6635 -4055
rect -6703 -4072 -6699 -4065
rect -6670 -4072 -6666 -4065
rect -6647 -4066 -6620 -4065
rect -6647 -4070 -6646 -4066
rect -6642 -4070 -6625 -4066
rect -6621 -4070 -6620 -4066
rect -6647 -4071 -6620 -4070
rect -6711 -4073 -6684 -4072
rect -6711 -4077 -6710 -4073
rect -6706 -4077 -6689 -4073
rect -6685 -4077 -6684 -4073
rect -6711 -4078 -6684 -4077
rect -6678 -4073 -6651 -4072
rect -6678 -4077 -6677 -4073
rect -6673 -4077 -6656 -4073
rect -6652 -4077 -6651 -4073
rect -6678 -4078 -6651 -4077
rect -6843 -4107 -6789 -4104
rect -6843 -4111 -6840 -4107
rect -6836 -4111 -6823 -4107
rect -6819 -4111 -6813 -4107
rect -6809 -4111 -6796 -4107
rect -6792 -4111 -6789 -4107
rect -6843 -4113 -6789 -4111
rect -6835 -4138 -6831 -4113
rect -6800 -4138 -6796 -4113
rect -6848 -4180 -6835 -4175
rect -6827 -4178 -6823 -4158
rect -6808 -4178 -6804 -4158
rect -6796 -4174 -6789 -4170
rect -6848 -4185 -6843 -4180
rect -6827 -4182 -6804 -4178
rect -6794 -4182 -6789 -4174
rect -6781 -4177 -6754 -4174
rect -6781 -4181 -6778 -4177
rect -6774 -4181 -6761 -4177
rect -6757 -4181 -6754 -4177
rect -6848 -4190 -6817 -4185
rect -6848 -4202 -6843 -4190
rect -6882 -4207 -6843 -4202
rect -6808 -4202 -6804 -4182
rect -6781 -4183 -6754 -4181
rect -6773 -4188 -6769 -4183
rect -6808 -4208 -6785 -4202
rect -6808 -4212 -6804 -4208
rect -6816 -4238 -6812 -4232
rect -6791 -4238 -6785 -4208
rect -6613 -4195 -6608 -4042
rect -6562 -4155 -6535 -4152
rect -6562 -4159 -6559 -4155
rect -6555 -4159 -6542 -4155
rect -6538 -4159 -6535 -4155
rect -6562 -4161 -6535 -4159
rect -6554 -4173 -6550 -4161
rect -6613 -4196 -6566 -4195
rect -6613 -4200 -6554 -4196
rect -6571 -4201 -6554 -4200
rect -6546 -4205 -6542 -4193
rect -6765 -4238 -6761 -4228
rect -6554 -4209 -6542 -4205
rect -6513 -4203 -6486 -4200
rect -6513 -4207 -6510 -4203
rect -6506 -4207 -6493 -4203
rect -6489 -4207 -6486 -4203
rect -6513 -4209 -6486 -4207
rect -6554 -4221 -6550 -4209
rect -6505 -4217 -6501 -4209
rect -6816 -4242 -6804 -4238
rect -7675 -4259 -7241 -4254
rect -7184 -4257 -6866 -4252
rect -6861 -4257 -6837 -4252
rect -6846 -4259 -6837 -4257
rect -6846 -4264 -6830 -4259
rect -6824 -4264 -6818 -4259
rect -6846 -4265 -6837 -4264
rect -6808 -4267 -6804 -4242
rect -6791 -4243 -6773 -4238
rect -6765 -4243 -6601 -4238
rect -6765 -4255 -6761 -4243
rect -6606 -4245 -6601 -4243
rect -6606 -4246 -6575 -4245
rect -6606 -4250 -6569 -4246
rect -6578 -4251 -6569 -4250
rect -6546 -4247 -6542 -4240
rect -6497 -4247 -6493 -4237
rect -6546 -4252 -6505 -4247
rect -6497 -4252 -6447 -4247
rect -6546 -4255 -6542 -4252
rect -6497 -4255 -6493 -4252
rect -7785 -4283 -7781 -4273
rect -7836 -4287 -7824 -4283
rect -8227 -4295 -8223 -4287
rect -8175 -4295 -8171 -4287
rect -8123 -4295 -8119 -4287
rect -8071 -4295 -8067 -4287
rect -8237 -4296 -8049 -4295
rect -8237 -4300 -8210 -4296
rect -8206 -4300 -8158 -4296
rect -8154 -4300 -8106 -4296
rect -8102 -4300 -8054 -4296
rect -8050 -4300 -8049 -4296
rect -8237 -4301 -8049 -4300
rect -7863 -4304 -7857 -4292
rect -7863 -4309 -7850 -4304
rect -7844 -4309 -7838 -4304
rect -8244 -4314 -8237 -4309
rect -8232 -4314 -8185 -4309
rect -8180 -4314 -8131 -4309
rect -8126 -4314 -8079 -4309
rect -7828 -4312 -7824 -4287
rect -7811 -4288 -7793 -4283
rect -7785 -4288 -6854 -4283
rect -7785 -4300 -7781 -4288
rect -7793 -4317 -7789 -4311
rect -7801 -4318 -7774 -4317
rect -7801 -4322 -7800 -4318
rect -7796 -4322 -7779 -4318
rect -7775 -4322 -7774 -4318
rect -7801 -4323 -7774 -4322
rect -6859 -4318 -6854 -4288
rect -6561 -4259 -6524 -4255
rect -6561 -4265 -6557 -4259
rect -6528 -4265 -6524 -4259
rect -6773 -4272 -6769 -4266
rect -6781 -4273 -6754 -4272
rect -6781 -4277 -6780 -4273
rect -6776 -4277 -6759 -4273
rect -6755 -4277 -6754 -4273
rect -6781 -4278 -6754 -4277
rect -6505 -4275 -6501 -4265
rect -6569 -4282 -6565 -4275
rect -6536 -4282 -6532 -4275
rect -6513 -4276 -6486 -4275
rect -6513 -4280 -6512 -4276
rect -6508 -4280 -6491 -4276
rect -6487 -4280 -6486 -4276
rect -6513 -4281 -6486 -4280
rect -6577 -4283 -6550 -4282
rect -6577 -4287 -6576 -4283
rect -6572 -4287 -6555 -4283
rect -6551 -4287 -6550 -4283
rect -6816 -4293 -6812 -4287
rect -6577 -4288 -6550 -4287
rect -6544 -4283 -6517 -4282
rect -6544 -4287 -6543 -4283
rect -6539 -4287 -6522 -4283
rect -6518 -4287 -6517 -4283
rect -6544 -4288 -6517 -4287
rect -6824 -4294 -6797 -4293
rect -6824 -4298 -6823 -4294
rect -6819 -4298 -6802 -4294
rect -6798 -4298 -6797 -4294
rect -6824 -4299 -6797 -4298
rect -6859 -4323 -6501 -4318
rect -7836 -4338 -7832 -4332
rect -7844 -4339 -7817 -4338
rect -7844 -4343 -7843 -4339
rect -7839 -4343 -7822 -4339
rect -7818 -4343 -7817 -4339
rect -7844 -4344 -7817 -4343
rect -6506 -4406 -6501 -4323
rect -6452 -4356 -6447 -4252
rect -6415 -4315 -6388 -4312
rect -6415 -4319 -6412 -4315
rect -6408 -4319 -6395 -4315
rect -6391 -4319 -6388 -4315
rect -6415 -4321 -6388 -4319
rect -6407 -4333 -6403 -4321
rect -6452 -4361 -6407 -4356
rect -6399 -4365 -6395 -4353
rect -6407 -4369 -6395 -4365
rect -6366 -4363 -6339 -4360
rect -6366 -4367 -6363 -4363
rect -6359 -4367 -6346 -4363
rect -6342 -4367 -6339 -4363
rect -6366 -4369 -6339 -4367
rect -6308 -4367 -6303 -3765
rect -6197 -4346 -6193 -4336
rect -5889 -4350 -5825 -4347
rect -5889 -4354 -5886 -4350
rect -5882 -4354 -5864 -4350
rect -5860 -4354 -5854 -4350
rect -5850 -4354 -5832 -4350
rect -5828 -4354 -5825 -4350
rect -6257 -4359 -6216 -4354
rect -6257 -4367 -6252 -4359
rect -6407 -4381 -6403 -4369
rect -6358 -4377 -6354 -4369
rect -6308 -4372 -6252 -4367
rect -6221 -4373 -6216 -4359
rect -6090 -4358 -5902 -4355
rect -5889 -4356 -5825 -4354
rect -6090 -4362 -6087 -4358
rect -6083 -4362 -6065 -4358
rect -6061 -4362 -6035 -4358
rect -6031 -4362 -6013 -4358
rect -6009 -4362 -5983 -4358
rect -5979 -4362 -5961 -4358
rect -5957 -4362 -5931 -4358
rect -5927 -4362 -5909 -4358
rect -5905 -4362 -5902 -4358
rect -6090 -4364 -5902 -4362
rect -5879 -4362 -5875 -4356
rect -5847 -4362 -5843 -4356
rect -6221 -4374 -6205 -4373
rect -6221 -4378 -6196 -4374
rect -6506 -4411 -6450 -4406
rect -6443 -4411 -6422 -4406
rect -6399 -4407 -6395 -4400
rect -6350 -4407 -6346 -4397
rect -6207 -4388 -6204 -4378
rect -6189 -4379 -6185 -4366
rect -6080 -4370 -6076 -4364
rect -6028 -4370 -6024 -4364
rect -5976 -4370 -5972 -4364
rect -5924 -4370 -5920 -4364
rect -6207 -4401 -6204 -4393
rect -6197 -4394 -6193 -4389
rect -6179 -4394 -6178 -4390
rect -6207 -4405 -6197 -4401
rect -6399 -4412 -6358 -4407
rect -6350 -4412 -6221 -4407
rect -5729 -4379 -5702 -4376
rect -5729 -4383 -5726 -4379
rect -5722 -4383 -5709 -4379
rect -5705 -4383 -5702 -4379
rect -5729 -4385 -5702 -4383
rect -6399 -4415 -6395 -4412
rect -6350 -4415 -6346 -4412
rect -6414 -4419 -6377 -4415
rect -6414 -4425 -6410 -4419
rect -6381 -4425 -6377 -4419
rect -6358 -4435 -6354 -4425
rect -6224 -4432 -6221 -4412
rect -6212 -4425 -6185 -4421
rect -6189 -4428 -6185 -4425
rect -6179 -4428 -6175 -4421
rect -6204 -4432 -6196 -4428
rect -6189 -4432 -6175 -4428
rect -6224 -4435 -6201 -4432
rect -6422 -4442 -6418 -4435
rect -6389 -4442 -6385 -4435
rect -6366 -4436 -6339 -4435
rect -6366 -4440 -6365 -4436
rect -6361 -4440 -6344 -4436
rect -6340 -4440 -6339 -4436
rect -6366 -4441 -6339 -4440
rect -6430 -4443 -6403 -4442
rect -6430 -4447 -6429 -4443
rect -6425 -4447 -6408 -4443
rect -6404 -4447 -6403 -4443
rect -6430 -4448 -6403 -4447
rect -6397 -4443 -6370 -4442
rect -6397 -4447 -6396 -4443
rect -6392 -4447 -6375 -4443
rect -6371 -4447 -6370 -4443
rect -6397 -4448 -6370 -4447
rect -6204 -4452 -6201 -4435
rect -6189 -4433 -6185 -4432
rect -6179 -4433 -6175 -4432
rect -6171 -4428 -6167 -4421
rect -6103 -4419 -6080 -4414
rect -6171 -4432 -6155 -4428
rect -6171 -4433 -6167 -4432
rect -6197 -4444 -6193 -4443
rect -6180 -4448 -6172 -4444
rect -6168 -4448 -6166 -4444
rect -6158 -4452 -6155 -4432
rect -6204 -4455 -6155 -4452
rect -6103 -4471 -6098 -4419
rect -6072 -4423 -6068 -4410
rect -6138 -4477 -6098 -4471
rect -6080 -4427 -6068 -4423
rect -6050 -4419 -6028 -4414
rect -6080 -4432 -6076 -4427
rect -6103 -4485 -6098 -4477
rect -6085 -4481 -6080 -4476
rect -6072 -4485 -6068 -4472
rect -6050 -4485 -6045 -4419
rect -6020 -4423 -6016 -4410
rect -5968 -4414 -5964 -4410
rect -5916 -4414 -5912 -4410
rect -5871 -4414 -5867 -4402
rect -5839 -4414 -5835 -4402
rect -5721 -4390 -5717 -4385
rect -6028 -4427 -6016 -4423
rect -5998 -4419 -5976 -4414
rect -5968 -4419 -5924 -4414
rect -5916 -4419 -5879 -4414
rect -5871 -4419 -5847 -4414
rect -5839 -4419 -5766 -4414
rect -6028 -4432 -6024 -4427
rect -6033 -4481 -6028 -4476
rect -6020 -4485 -6016 -4472
rect -5998 -4485 -5993 -4419
rect -5979 -4442 -5976 -4437
rect -5968 -4446 -5964 -4419
rect -5976 -4477 -5972 -4466
rect -5976 -4481 -5964 -4477
rect -6103 -4490 -6080 -4485
rect -6072 -4490 -6028 -4485
rect -6020 -4490 -5976 -4485
rect -6072 -4493 -6068 -4490
rect -6020 -4493 -6016 -4490
rect -5968 -4493 -5964 -4481
rect -5946 -4485 -5941 -4419
rect -5927 -4442 -5924 -4437
rect -5916 -4446 -5912 -4419
rect -5871 -4422 -5867 -4419
rect -5839 -4422 -5835 -4419
rect -5771 -4440 -5766 -4419
rect -5713 -4440 -5709 -4430
rect -5879 -4449 -5875 -4442
rect -5847 -4449 -5843 -4442
rect -5771 -4445 -5721 -4440
rect -5713 -4445 -5700 -4440
rect -5889 -4451 -5825 -4449
rect -5889 -4455 -5887 -4451
rect -5883 -4455 -5863 -4451
rect -5859 -4455 -5855 -4451
rect -5851 -4455 -5831 -4451
rect -5827 -4455 -5825 -4451
rect -5889 -4457 -5825 -4455
rect -5713 -4457 -5709 -4445
rect -5924 -4477 -5920 -4466
rect -5721 -4474 -5717 -4468
rect -5729 -4475 -5702 -4474
rect -5924 -4481 -5912 -4477
rect -5729 -4479 -5728 -4475
rect -5724 -4479 -5707 -4475
rect -5703 -4479 -5702 -4475
rect -5729 -4480 -5702 -4479
rect -5946 -4490 -5924 -4485
rect -5916 -4493 -5912 -4481
rect -6080 -4521 -6076 -4513
rect -6028 -4521 -6024 -4513
rect -5976 -4521 -5972 -4513
rect -5924 -4521 -5920 -4513
rect -6090 -4522 -5902 -4521
rect -6090 -4526 -6063 -4522
rect -6059 -4526 -6011 -4522
rect -6007 -4526 -5959 -4522
rect -5955 -4526 -5907 -4522
rect -5903 -4526 -5902 -4522
rect -6090 -4527 -5902 -4526
rect -6097 -4540 -6090 -4535
rect -6085 -4540 -6038 -4535
rect -6033 -4540 -5984 -4535
rect -5979 -4540 -5932 -4535
rect -7609 -4664 -7555 -4661
rect -7736 -4670 -7709 -4667
rect -7609 -4668 -7606 -4664
rect -7602 -4668 -7589 -4664
rect -7585 -4668 -7579 -4664
rect -7575 -4668 -7562 -4664
rect -7558 -4668 -7555 -4664
rect -7609 -4670 -7555 -4668
rect -7911 -4677 -7841 -4672
rect -7736 -4674 -7733 -4670
rect -7729 -4674 -7716 -4670
rect -7712 -4674 -7709 -4670
rect -7736 -4676 -7709 -4674
rect -8047 -4687 -7983 -4684
rect -8047 -4691 -8044 -4687
rect -8040 -4691 -8022 -4687
rect -8018 -4691 -8012 -4687
rect -8008 -4691 -7990 -4687
rect -7986 -4691 -7983 -4687
rect -8248 -4695 -8060 -4692
rect -8047 -4693 -7983 -4691
rect -8248 -4699 -8245 -4695
rect -8241 -4699 -8223 -4695
rect -8219 -4699 -8193 -4695
rect -8189 -4699 -8171 -4695
rect -8167 -4699 -8141 -4695
rect -8137 -4699 -8119 -4695
rect -8115 -4699 -8089 -4695
rect -8085 -4699 -8067 -4695
rect -8063 -4699 -8060 -4695
rect -8248 -4701 -8060 -4699
rect -8037 -4699 -8033 -4693
rect -8005 -4699 -8001 -4693
rect -8238 -4707 -8234 -4701
rect -8186 -4707 -8182 -4701
rect -8134 -4707 -8130 -4701
rect -8082 -4707 -8078 -4701
rect -8261 -4756 -8238 -4751
rect -8261 -4822 -8256 -4756
rect -8230 -4760 -8226 -4747
rect -8238 -4764 -8226 -4760
rect -8208 -4756 -8186 -4751
rect -8238 -4769 -8234 -4764
rect -8243 -4818 -8238 -4813
rect -8230 -4822 -8226 -4809
rect -8208 -4822 -8203 -4756
rect -8178 -4760 -8174 -4747
rect -8126 -4751 -8122 -4747
rect -8074 -4751 -8070 -4747
rect -8029 -4751 -8025 -4739
rect -7997 -4751 -7993 -4739
rect -7911 -4751 -7906 -4677
rect -7876 -4681 -7870 -4680
rect -7876 -4685 -7875 -4681
rect -7871 -4685 -7870 -4681
rect -7876 -4688 -7870 -4685
rect -7841 -4688 -7836 -4677
rect -7791 -4683 -7782 -4680
rect -7791 -4687 -7789 -4683
rect -7785 -4687 -7782 -4683
rect -7791 -4688 -7782 -4687
rect -7876 -4692 -7864 -4688
rect -7876 -4702 -7870 -4692
rect -7806 -4692 -7782 -4688
rect -7728 -4684 -7724 -4676
rect -7841 -4700 -7826 -4696
rect -7791 -4700 -7782 -4692
rect -7756 -4696 -7743 -4692
rect -7756 -4699 -7752 -4696
rect -7876 -4706 -7875 -4702
rect -7871 -4706 -7870 -4702
rect -7876 -4707 -7870 -4706
rect -7841 -4710 -7836 -4700
rect -7791 -4704 -7789 -4700
rect -7785 -4704 -7782 -4700
rect -7791 -4707 -7782 -4704
rect -7764 -4710 -7760 -4707
rect -7812 -4714 -7760 -4710
rect -7812 -4719 -7808 -4714
rect -7871 -4724 -7808 -4719
rect -8186 -4764 -8174 -4760
rect -8156 -4756 -8134 -4751
rect -8126 -4756 -8082 -4751
rect -8074 -4756 -8037 -4751
rect -8029 -4756 -8005 -4751
rect -7997 -4756 -7906 -4751
rect -8186 -4769 -8182 -4764
rect -8191 -4818 -8186 -4813
rect -8178 -4822 -8174 -4809
rect -8156 -4822 -8151 -4756
rect -8137 -4779 -8134 -4774
rect -8126 -4783 -8122 -4756
rect -8134 -4814 -8130 -4803
rect -8134 -4818 -8122 -4814
rect -8261 -4827 -8238 -4822
rect -8230 -4827 -8186 -4822
rect -8178 -4827 -8134 -4822
rect -8230 -4830 -8226 -4827
rect -8178 -4830 -8174 -4827
rect -8126 -4830 -8122 -4818
rect -8104 -4822 -8099 -4756
rect -8085 -4779 -8082 -4774
rect -8074 -4783 -8070 -4756
rect -8029 -4759 -8025 -4756
rect -7997 -4759 -7993 -4756
rect -8037 -4786 -8033 -4779
rect -8005 -4786 -8001 -4779
rect -8047 -4788 -7983 -4786
rect -8047 -4792 -8045 -4788
rect -8041 -4792 -8021 -4788
rect -8017 -4792 -8013 -4788
rect -8009 -4792 -7989 -4788
rect -7985 -4792 -7983 -4788
rect -8047 -4794 -7983 -4792
rect -8082 -4814 -8078 -4803
rect -8082 -4818 -8070 -4814
rect -8104 -4827 -8082 -4822
rect -8074 -4830 -8070 -4818
rect -8238 -4858 -8234 -4850
rect -8186 -4858 -8182 -4850
rect -8134 -4858 -8130 -4850
rect -8082 -4858 -8078 -4850
rect -8248 -4859 -8060 -4858
rect -8248 -4863 -8221 -4859
rect -8217 -4863 -8169 -4859
rect -8165 -4863 -8117 -4859
rect -8113 -4863 -8065 -4859
rect -8061 -4863 -8060 -4859
rect -8248 -4864 -8060 -4863
rect -8255 -4877 -8248 -4872
rect -8243 -4877 -8196 -4872
rect -8191 -4877 -8142 -4872
rect -8137 -4877 -8090 -4872
rect -8034 -4999 -7970 -4996
rect -8034 -5003 -8031 -4999
rect -8027 -5003 -8009 -4999
rect -8005 -5003 -7999 -4999
rect -7995 -5003 -7977 -4999
rect -7973 -5003 -7970 -4999
rect -8235 -5007 -8047 -5004
rect -8034 -5005 -7970 -5003
rect -8235 -5011 -8232 -5007
rect -8228 -5011 -8210 -5007
rect -8206 -5011 -8180 -5007
rect -8176 -5011 -8158 -5007
rect -8154 -5011 -8128 -5007
rect -8124 -5011 -8106 -5007
rect -8102 -5011 -8076 -5007
rect -8072 -5011 -8054 -5007
rect -8050 -5011 -8047 -5007
rect -8235 -5013 -8047 -5011
rect -8024 -5011 -8020 -5005
rect -7992 -5011 -7988 -5005
rect -8225 -5019 -8221 -5013
rect -8173 -5019 -8169 -5013
rect -8121 -5019 -8117 -5013
rect -8069 -5019 -8065 -5013
rect -8248 -5068 -8225 -5063
rect -8248 -5134 -8243 -5068
rect -8217 -5072 -8213 -5059
rect -8225 -5076 -8213 -5072
rect -8195 -5068 -8173 -5063
rect -8225 -5081 -8221 -5076
rect -8230 -5130 -8225 -5125
rect -8217 -5134 -8213 -5121
rect -8195 -5134 -8190 -5068
rect -8165 -5072 -8161 -5059
rect -8113 -5063 -8109 -5059
rect -8061 -5063 -8057 -5059
rect -8016 -5063 -8012 -5051
rect -7984 -5063 -7980 -5051
rect -8173 -5076 -8161 -5072
rect -8143 -5068 -8121 -5063
rect -8113 -5068 -8069 -5063
rect -8061 -5068 -8024 -5063
rect -8016 -5068 -7992 -5063
rect -7984 -5068 -7976 -5063
rect -8173 -5081 -8169 -5076
rect -8178 -5130 -8173 -5125
rect -8165 -5134 -8161 -5121
rect -8143 -5134 -8138 -5068
rect -8124 -5091 -8121 -5086
rect -8113 -5095 -8109 -5068
rect -8121 -5126 -8117 -5115
rect -8121 -5130 -8109 -5126
rect -8248 -5139 -8225 -5134
rect -8217 -5139 -8173 -5134
rect -8165 -5139 -8121 -5134
rect -8217 -5142 -8213 -5139
rect -8165 -5142 -8161 -5139
rect -8113 -5142 -8109 -5130
rect -8091 -5134 -8086 -5068
rect -8072 -5091 -8069 -5086
rect -8061 -5095 -8057 -5068
rect -8016 -5071 -8012 -5068
rect -7984 -5071 -7980 -5068
rect -8024 -5098 -8020 -5091
rect -7992 -5098 -7988 -5091
rect -7911 -5097 -7906 -4756
rect -7876 -4732 -7870 -4731
rect -7876 -4736 -7875 -4732
rect -7871 -4736 -7870 -4732
rect -7876 -4739 -7870 -4736
rect -7841 -4739 -7836 -4724
rect -7756 -4730 -7752 -4707
rect -7749 -4714 -7743 -4696
rect -7720 -4714 -7716 -4704
rect -7601 -4695 -7597 -4670
rect -7566 -4695 -7562 -4670
rect -7749 -4719 -7728 -4714
rect -7720 -4719 -7658 -4714
rect -7720 -4722 -7716 -4719
rect -7791 -4734 -7782 -4731
rect -7791 -4738 -7789 -4734
rect -7785 -4738 -7782 -4734
rect -7791 -4739 -7782 -4738
rect -7876 -4743 -7864 -4739
rect -7876 -4753 -7870 -4743
rect -7806 -4743 -7782 -4739
rect -7841 -4751 -7826 -4747
rect -7791 -4751 -7782 -4743
rect -7876 -4757 -7875 -4753
rect -7871 -4757 -7870 -4753
rect -7876 -4758 -7870 -4757
rect -7841 -4762 -7836 -4751
rect -7791 -4755 -7789 -4751
rect -7785 -4755 -7782 -4751
rect -7791 -4758 -7782 -4755
rect -7764 -4762 -7760 -4740
rect -7728 -4742 -7724 -4732
rect -7736 -4743 -7709 -4742
rect -7736 -4747 -7735 -4743
rect -7731 -4747 -7714 -4743
rect -7710 -4747 -7709 -4743
rect -7736 -4748 -7709 -4747
rect -7841 -4765 -7760 -4762
rect -7869 -5001 -7815 -4998
rect -7869 -5005 -7866 -5001
rect -7862 -5005 -7849 -5001
rect -7845 -5005 -7839 -5001
rect -7835 -5005 -7822 -5001
rect -7818 -5005 -7815 -5001
rect -7869 -5007 -7815 -5005
rect -7861 -5032 -7857 -5007
rect -7826 -5032 -7822 -5007
rect -7874 -5074 -7861 -5069
rect -7853 -5072 -7849 -5052
rect -7834 -5072 -7830 -5052
rect -7822 -5068 -7815 -5064
rect -7874 -5079 -7869 -5074
rect -7853 -5076 -7830 -5072
rect -7820 -5076 -7815 -5068
rect -7807 -5071 -7780 -5068
rect -7807 -5075 -7804 -5071
rect -7800 -5075 -7787 -5071
rect -7783 -5075 -7780 -5071
rect -7874 -5084 -7843 -5079
rect -7874 -5097 -7869 -5084
rect -8034 -5100 -7970 -5098
rect -8034 -5104 -8032 -5100
rect -8028 -5104 -8008 -5100
rect -8004 -5104 -8000 -5100
rect -7996 -5104 -7976 -5100
rect -7972 -5104 -7970 -5100
rect -7911 -5102 -7869 -5097
rect -7834 -5096 -7830 -5076
rect -7807 -5077 -7780 -5075
rect -7799 -5082 -7795 -5077
rect -7834 -5102 -7811 -5096
rect -8034 -5106 -7970 -5104
rect -7834 -5106 -7830 -5102
rect -8069 -5126 -8065 -5115
rect -8069 -5130 -8057 -5126
rect -8091 -5139 -8069 -5134
rect -8061 -5142 -8057 -5130
rect -7842 -5132 -7838 -5126
rect -7817 -5132 -7811 -5102
rect -7690 -5114 -7685 -4719
rect -7663 -4759 -7658 -4719
rect -7614 -4737 -7601 -4732
rect -7593 -4735 -7589 -4715
rect -7574 -4735 -7570 -4715
rect -7562 -4731 -7555 -4727
rect -7614 -4742 -7609 -4737
rect -7593 -4739 -7570 -4735
rect -7560 -4739 -7555 -4731
rect -7547 -4734 -7520 -4731
rect -7547 -4738 -7544 -4734
rect -7540 -4738 -7527 -4734
rect -7523 -4738 -7520 -4734
rect -7614 -4747 -7583 -4742
rect -7614 -4759 -7609 -4747
rect -7663 -4764 -7637 -4759
rect -7632 -4764 -7628 -4759
rect -7623 -4764 -7609 -4759
rect -7574 -4759 -7570 -4739
rect -7547 -4740 -7520 -4738
rect -7539 -4745 -7535 -4740
rect -7574 -4765 -7551 -4759
rect -7574 -4769 -7570 -4765
rect -7582 -4795 -7578 -4789
rect -7557 -4795 -7551 -4765
rect -7531 -4795 -7527 -4785
rect -7651 -4805 -7603 -4798
rect -7582 -4799 -7570 -4795
rect -7610 -4816 -7603 -4805
rect -7610 -4821 -7596 -4816
rect -7590 -4821 -7584 -4816
rect -7574 -4824 -7570 -4799
rect -7557 -4800 -7539 -4795
rect -7531 -4800 -7464 -4795
rect -7531 -4812 -7527 -4800
rect -7539 -4829 -7535 -4823
rect -7547 -4830 -7520 -4829
rect -7547 -4834 -7546 -4830
rect -7542 -4834 -7525 -4830
rect -7521 -4834 -7520 -4830
rect -7547 -4835 -7520 -4834
rect -7582 -4850 -7578 -4844
rect -7469 -4846 -7464 -4800
rect -7443 -4805 -7416 -4802
rect -7443 -4809 -7440 -4805
rect -7436 -4809 -7423 -4805
rect -7419 -4809 -7416 -4805
rect -7443 -4811 -7416 -4809
rect -7435 -4823 -7431 -4811
rect -7590 -4851 -7563 -4850
rect -7469 -4851 -7435 -4846
rect -7590 -4855 -7589 -4851
rect -7585 -4855 -7568 -4851
rect -7564 -4855 -7563 -4851
rect -7427 -4855 -7423 -4843
rect -7590 -4856 -7563 -4855
rect -7435 -4859 -7423 -4855
rect -7394 -4853 -7367 -4850
rect -7394 -4857 -7391 -4853
rect -7387 -4857 -7374 -4853
rect -7370 -4857 -7367 -4853
rect -7394 -4859 -7367 -4857
rect -7608 -4869 -7554 -4866
rect -7608 -4873 -7605 -4869
rect -7601 -4873 -7588 -4869
rect -7584 -4873 -7578 -4869
rect -7574 -4873 -7561 -4869
rect -7557 -4873 -7554 -4869
rect -7608 -4875 -7554 -4873
rect -7435 -4871 -7431 -4859
rect -7386 -4867 -7382 -4859
rect -7600 -4900 -7596 -4875
rect -7565 -4900 -7561 -4875
rect -7613 -4942 -7600 -4937
rect -7592 -4940 -7588 -4920
rect -7487 -4895 -7459 -4894
rect -7487 -4896 -7458 -4895
rect -7487 -4899 -7450 -4896
rect -7573 -4940 -7569 -4920
rect -7561 -4936 -7554 -4932
rect -7613 -4947 -7608 -4942
rect -7592 -4944 -7569 -4940
rect -7559 -4944 -7554 -4936
rect -7546 -4939 -7519 -4936
rect -7546 -4943 -7543 -4939
rect -7539 -4943 -7526 -4939
rect -7522 -4943 -7519 -4939
rect -7613 -4952 -7582 -4947
rect -7613 -4963 -7608 -4952
rect -7616 -4968 -7608 -4963
rect -7573 -4964 -7569 -4944
rect -7546 -4945 -7519 -4943
rect -7538 -4950 -7534 -4945
rect -7573 -4970 -7550 -4964
rect -7573 -4974 -7569 -4970
rect -7581 -5000 -7577 -4994
rect -7556 -5000 -7550 -4970
rect -7530 -5000 -7526 -4990
rect -7487 -5000 -7482 -4899
rect -7464 -4901 -7450 -4899
rect -7427 -4897 -7423 -4890
rect -7378 -4897 -7374 -4887
rect -7427 -4902 -7386 -4897
rect -7378 -4902 -7338 -4897
rect -7427 -4905 -7423 -4902
rect -7378 -4905 -7374 -4902
rect -7442 -4909 -7405 -4905
rect -7442 -4915 -7438 -4909
rect -7409 -4915 -7405 -4909
rect -7386 -4925 -7382 -4915
rect -7450 -4932 -7446 -4925
rect -7417 -4932 -7413 -4925
rect -7394 -4926 -7367 -4925
rect -7394 -4930 -7393 -4926
rect -7389 -4930 -7372 -4926
rect -7368 -4930 -7367 -4926
rect -7394 -4931 -7367 -4930
rect -7458 -4933 -7431 -4932
rect -7458 -4937 -7457 -4933
rect -7453 -4937 -7436 -4933
rect -7432 -4937 -7431 -4933
rect -7458 -4938 -7431 -4937
rect -7425 -4933 -7398 -4932
rect -7425 -4937 -7424 -4933
rect -7420 -4937 -7403 -4933
rect -7399 -4937 -7398 -4933
rect -7425 -4938 -7398 -4937
rect -7343 -4959 -7338 -4902
rect -7297 -4918 -7270 -4915
rect -7297 -4922 -7294 -4918
rect -7290 -4922 -7277 -4918
rect -7273 -4922 -7270 -4918
rect -7297 -4924 -7270 -4922
rect -7289 -4936 -7285 -4924
rect -7343 -4964 -7289 -4959
rect -7281 -4968 -7277 -4956
rect -7115 -4957 -7111 -4947
rect -6808 -4959 -6744 -4956
rect -6808 -4963 -6805 -4959
rect -6801 -4963 -6783 -4959
rect -6779 -4963 -6773 -4959
rect -6769 -4963 -6751 -4959
rect -6747 -4963 -6744 -4959
rect -7581 -5004 -7569 -5000
rect -7602 -5026 -7595 -5021
rect -7589 -5026 -7583 -5021
rect -7573 -5029 -7569 -5004
rect -7556 -5005 -7538 -5000
rect -7530 -5005 -7482 -5000
rect -7289 -4972 -7277 -4968
rect -7248 -4966 -7221 -4963
rect -7248 -4970 -7245 -4966
rect -7241 -4970 -7228 -4966
rect -7224 -4970 -7221 -4966
rect -7248 -4972 -7221 -4970
rect -7009 -4967 -6821 -4964
rect -6808 -4965 -6744 -4963
rect -7009 -4971 -7006 -4967
rect -7002 -4971 -6984 -4967
rect -6980 -4971 -6954 -4967
rect -6950 -4971 -6932 -4967
rect -6928 -4971 -6902 -4967
rect -6898 -4971 -6880 -4967
rect -6876 -4971 -6850 -4967
rect -6846 -4971 -6828 -4967
rect -6824 -4971 -6821 -4967
rect -7289 -4984 -7285 -4972
rect -7240 -4980 -7236 -4972
rect -7009 -4973 -6821 -4971
rect -6798 -4971 -6794 -4965
rect -6766 -4971 -6762 -4965
rect -7530 -5017 -7526 -5005
rect -7313 -5010 -7304 -5009
rect -7357 -5015 -7331 -5010
rect -7321 -5014 -7304 -5010
rect -7281 -5010 -7277 -5003
rect -7232 -5010 -7228 -5000
rect -7120 -4989 -7114 -4985
rect -7107 -4990 -7103 -4977
rect -6999 -4979 -6995 -4973
rect -6947 -4979 -6943 -4973
rect -6895 -4979 -6891 -4973
rect -6843 -4979 -6839 -4973
rect -7125 -4999 -7122 -4990
rect -7321 -5015 -7310 -5014
rect -7281 -5015 -7240 -5010
rect -7232 -5015 -7144 -5010
rect -7538 -5034 -7534 -5028
rect -7546 -5035 -7519 -5034
rect -7546 -5039 -7545 -5035
rect -7541 -5039 -7524 -5035
rect -7520 -5039 -7519 -5035
rect -7546 -5040 -7519 -5039
rect -7581 -5055 -7577 -5049
rect -7589 -5056 -7562 -5055
rect -7589 -5060 -7588 -5056
rect -7584 -5060 -7567 -5056
rect -7563 -5060 -7562 -5056
rect -7589 -5061 -7562 -5060
rect -7791 -5132 -7787 -5122
rect -7357 -5132 -7352 -5015
rect -7281 -5018 -7277 -5015
rect -7232 -5018 -7228 -5015
rect -7296 -5022 -7259 -5018
rect -7296 -5028 -7292 -5022
rect -7263 -5028 -7259 -5022
rect -7240 -5038 -7236 -5028
rect -7304 -5045 -7300 -5038
rect -7271 -5045 -7267 -5038
rect -7248 -5039 -7221 -5038
rect -7248 -5043 -7247 -5039
rect -7243 -5043 -7226 -5039
rect -7222 -5043 -7221 -5039
rect -7248 -5044 -7221 -5043
rect -7149 -5042 -7144 -5015
rect -7125 -5012 -7122 -5004
rect -7115 -5005 -7111 -5000
rect -7097 -5005 -7096 -5001
rect -7125 -5016 -7115 -5012
rect -6695 -4999 -6668 -4996
rect -6695 -5003 -6692 -4999
rect -6688 -5003 -6675 -4999
rect -6671 -5003 -6668 -4999
rect -6695 -5005 -6668 -5003
rect -7022 -5028 -6999 -5023
rect -7129 -5036 -7103 -5032
rect -7107 -5039 -7103 -5036
rect -7097 -5039 -7093 -5032
rect -7122 -5042 -7114 -5039
rect -7149 -5043 -7114 -5042
rect -7107 -5043 -7093 -5039
rect -7312 -5046 -7285 -5045
rect -7312 -5050 -7311 -5046
rect -7307 -5050 -7290 -5046
rect -7286 -5050 -7285 -5046
rect -7312 -5051 -7285 -5050
rect -7279 -5046 -7252 -5045
rect -7149 -5046 -7119 -5043
rect -7279 -5050 -7278 -5046
rect -7274 -5050 -7257 -5046
rect -7253 -5050 -7252 -5046
rect -7279 -5051 -7252 -5050
rect -7122 -5063 -7119 -5046
rect -7107 -5044 -7103 -5043
rect -7097 -5044 -7093 -5043
rect -7089 -5039 -7085 -5032
rect -7089 -5043 -7073 -5039
rect -7089 -5044 -7085 -5043
rect -7115 -5055 -7111 -5054
rect -7098 -5059 -7090 -5055
rect -7086 -5059 -7084 -5055
rect -7076 -5063 -7073 -5043
rect -7122 -5066 -7073 -5063
rect -7022 -5089 -7017 -5028
rect -6991 -5032 -6987 -5019
rect -6999 -5036 -6987 -5032
rect -6969 -5028 -6947 -5023
rect -6999 -5041 -6995 -5036
rect -7062 -5094 -7017 -5089
rect -7004 -5090 -6999 -5085
rect -6991 -5094 -6987 -5081
rect -6969 -5094 -6964 -5028
rect -6939 -5032 -6935 -5019
rect -6887 -5023 -6883 -5019
rect -6835 -5023 -6831 -5019
rect -6790 -5023 -6786 -5011
rect -6758 -5023 -6754 -5011
rect -6687 -5010 -6683 -5005
rect -6947 -5036 -6935 -5032
rect -6917 -5028 -6895 -5023
rect -6887 -5028 -6843 -5023
rect -6835 -5028 -6798 -5023
rect -6790 -5028 -6766 -5023
rect -6758 -5028 -6713 -5023
rect -6947 -5041 -6943 -5036
rect -6952 -5090 -6947 -5085
rect -6939 -5094 -6935 -5081
rect -6917 -5094 -6912 -5028
rect -6898 -5051 -6895 -5046
rect -6887 -5055 -6883 -5028
rect -6895 -5086 -6891 -5075
rect -6895 -5090 -6883 -5086
rect -7022 -5099 -6999 -5094
rect -6991 -5099 -6947 -5094
rect -6939 -5099 -6895 -5094
rect -6991 -5102 -6987 -5099
rect -6939 -5102 -6935 -5099
rect -6887 -5102 -6883 -5090
rect -6865 -5094 -6860 -5028
rect -6846 -5051 -6843 -5046
rect -6835 -5055 -6831 -5028
rect -6790 -5031 -6786 -5028
rect -6758 -5031 -6754 -5028
rect -6798 -5058 -6794 -5051
rect -6766 -5058 -6762 -5051
rect -6808 -5060 -6744 -5058
rect -6808 -5064 -6806 -5060
rect -6802 -5064 -6782 -5060
rect -6778 -5064 -6774 -5060
rect -6770 -5064 -6750 -5060
rect -6746 -5064 -6744 -5060
rect -6808 -5066 -6744 -5064
rect -6718 -5061 -6713 -5028
rect -6679 -5060 -6675 -5050
rect -3990 -5057 -3986 -5047
rect -6697 -5061 -6687 -5060
rect -6718 -5065 -6687 -5061
rect -6679 -5065 -6666 -5060
rect -6718 -5066 -6691 -5065
rect -6843 -5086 -6839 -5075
rect -6679 -5077 -6675 -5065
rect -6843 -5090 -6831 -5086
rect -6865 -5099 -6843 -5094
rect -6835 -5102 -6831 -5090
rect -6687 -5094 -6683 -5088
rect -4000 -5089 -3989 -5085
rect -6695 -5095 -6668 -5094
rect -6695 -5099 -6694 -5095
rect -6690 -5099 -6673 -5095
rect -6669 -5099 -6668 -5095
rect -6695 -5100 -6668 -5099
rect -4000 -5099 -3997 -5089
rect -3982 -5090 -3978 -5077
rect -4000 -5112 -3997 -5104
rect -3990 -5105 -3986 -5100
rect -3972 -5105 -3971 -5101
rect -4000 -5116 -3990 -5112
rect -6999 -5130 -6995 -5122
rect -6947 -5130 -6943 -5122
rect -6895 -5130 -6891 -5122
rect -6843 -5130 -6839 -5122
rect -7842 -5136 -7830 -5132
rect -7869 -5153 -7863 -5143
rect -7869 -5158 -7856 -5153
rect -7850 -5158 -7844 -5153
rect -7834 -5161 -7830 -5136
rect -7817 -5137 -7799 -5132
rect -7791 -5137 -7352 -5132
rect -7009 -5131 -6821 -5130
rect -7009 -5135 -6982 -5131
rect -6978 -5135 -6930 -5131
rect -6926 -5135 -6878 -5131
rect -6874 -5135 -6826 -5131
rect -6822 -5135 -6821 -5131
rect -7009 -5136 -6821 -5135
rect -7791 -5149 -7787 -5137
rect -3982 -5139 -3978 -5132
rect -3972 -5139 -3968 -5132
rect -3997 -5143 -3989 -5139
rect -3982 -5143 -3968 -5139
rect -8225 -5170 -8221 -5162
rect -8173 -5170 -8169 -5162
rect -8121 -5170 -8117 -5162
rect -8069 -5170 -8065 -5162
rect -8235 -5171 -8047 -5170
rect -8235 -5175 -8208 -5171
rect -8204 -5175 -8156 -5171
rect -8152 -5175 -8104 -5171
rect -8100 -5175 -8052 -5171
rect -8048 -5175 -8047 -5171
rect -8235 -5176 -8047 -5175
rect -7016 -5149 -7009 -5144
rect -7004 -5149 -6957 -5144
rect -6952 -5149 -6903 -5144
rect -6898 -5149 -6851 -5144
rect -7690 -5157 -7685 -5153
rect -7799 -5166 -7795 -5160
rect -7807 -5167 -7780 -5166
rect -7807 -5171 -7806 -5167
rect -7802 -5171 -7785 -5167
rect -7781 -5171 -7780 -5167
rect -7807 -5172 -7780 -5171
rect -8242 -5189 -8235 -5184
rect -8230 -5189 -8183 -5184
rect -8178 -5189 -8129 -5184
rect -8124 -5189 -8077 -5184
rect -7842 -5187 -7838 -5181
rect -7850 -5188 -7823 -5187
rect -7850 -5192 -7849 -5188
rect -7845 -5192 -7828 -5188
rect -7824 -5192 -7823 -5188
rect -7850 -5193 -7823 -5192
rect -7689 -5207 -7685 -5157
rect -3997 -5163 -3994 -5143
rect -3982 -5144 -3978 -5143
rect -3972 -5144 -3968 -5143
rect -3964 -5139 -3960 -5132
rect -3964 -5143 -3948 -5139
rect -3964 -5144 -3960 -5143
rect -3990 -5155 -3986 -5154
rect -3973 -5159 -3965 -5155
rect -3961 -5159 -3959 -5155
rect -3951 -5163 -3948 -5143
rect -3997 -5166 -3948 -5163
rect -7689 -5211 -7427 -5207
rect -7652 -5302 -7584 -5295
rect -8047 -5393 -7983 -5390
rect -8047 -5397 -8044 -5393
rect -8040 -5397 -8022 -5393
rect -8018 -5397 -8012 -5393
rect -8008 -5397 -7990 -5393
rect -7986 -5397 -7983 -5393
rect -8248 -5401 -8060 -5398
rect -8047 -5399 -7983 -5397
rect -8248 -5405 -8245 -5401
rect -8241 -5405 -8223 -5401
rect -8219 -5405 -8193 -5401
rect -8189 -5405 -8171 -5401
rect -8167 -5405 -8141 -5401
rect -8137 -5405 -8119 -5401
rect -8115 -5405 -8089 -5401
rect -8085 -5405 -8067 -5401
rect -8063 -5405 -8060 -5401
rect -8248 -5407 -8060 -5405
rect -8037 -5405 -8033 -5399
rect -8005 -5405 -8001 -5399
rect -8238 -5413 -8234 -5407
rect -8186 -5413 -8182 -5407
rect -8134 -5413 -8130 -5407
rect -8082 -5413 -8078 -5407
rect -7758 -5432 -7731 -5429
rect -8261 -5462 -8238 -5457
rect -8261 -5528 -8256 -5462
rect -8230 -5466 -8226 -5453
rect -8238 -5470 -8226 -5466
rect -8208 -5462 -8186 -5457
rect -8238 -5475 -8234 -5470
rect -8243 -5524 -8238 -5519
rect -8230 -5528 -8226 -5515
rect -8208 -5528 -8203 -5462
rect -8178 -5466 -8174 -5453
rect -8126 -5457 -8122 -5453
rect -8074 -5457 -8070 -5453
rect -8029 -5457 -8025 -5445
rect -7997 -5457 -7993 -5445
rect -7929 -5439 -7863 -5434
rect -7758 -5436 -7755 -5432
rect -7751 -5436 -7738 -5432
rect -7734 -5436 -7731 -5432
rect -7758 -5438 -7731 -5436
rect -7929 -5457 -7924 -5439
rect -8186 -5470 -8174 -5466
rect -8156 -5462 -8134 -5457
rect -8126 -5462 -8082 -5457
rect -8074 -5462 -8037 -5457
rect -8029 -5462 -8005 -5457
rect -7997 -5462 -7924 -5457
rect -8186 -5475 -8182 -5470
rect -8191 -5524 -8186 -5519
rect -8178 -5528 -8174 -5515
rect -8156 -5528 -8151 -5462
rect -8137 -5485 -8134 -5480
rect -8126 -5489 -8122 -5462
rect -8134 -5520 -8130 -5509
rect -8134 -5524 -8122 -5520
rect -8261 -5533 -8238 -5528
rect -8230 -5533 -8186 -5528
rect -8178 -5533 -8134 -5528
rect -8230 -5536 -8226 -5533
rect -8178 -5536 -8174 -5533
rect -8126 -5536 -8122 -5524
rect -8104 -5528 -8099 -5462
rect -8085 -5485 -8082 -5480
rect -8074 -5489 -8070 -5462
rect -8029 -5465 -8025 -5462
rect -7997 -5465 -7993 -5462
rect -8037 -5492 -8033 -5485
rect -8005 -5492 -8001 -5485
rect -8047 -5494 -7983 -5492
rect -8047 -5498 -8045 -5494
rect -8041 -5498 -8021 -5494
rect -8017 -5498 -8013 -5494
rect -8009 -5498 -7989 -5494
rect -7985 -5498 -7983 -5494
rect -8047 -5500 -7983 -5498
rect -8082 -5520 -8078 -5509
rect -8082 -5524 -8070 -5520
rect -8104 -5533 -8082 -5528
rect -8074 -5536 -8070 -5524
rect -8238 -5564 -8234 -5556
rect -8186 -5564 -8182 -5556
rect -8134 -5564 -8130 -5556
rect -8082 -5564 -8078 -5556
rect -8248 -5565 -8060 -5564
rect -8248 -5569 -8221 -5565
rect -8217 -5569 -8169 -5565
rect -8165 -5569 -8117 -5565
rect -8113 -5569 -8065 -5565
rect -8061 -5569 -8060 -5565
rect -8248 -5570 -8060 -5569
rect -8255 -5583 -8248 -5578
rect -8243 -5583 -8196 -5578
rect -8191 -5583 -8142 -5578
rect -8137 -5583 -8090 -5578
rect -8044 -5642 -7980 -5639
rect -8044 -5646 -8041 -5642
rect -8037 -5646 -8019 -5642
rect -8015 -5646 -8009 -5642
rect -8005 -5646 -7987 -5642
rect -7983 -5646 -7980 -5642
rect -8245 -5650 -8057 -5647
rect -8044 -5648 -7980 -5646
rect -8245 -5654 -8242 -5650
rect -8238 -5654 -8220 -5650
rect -8216 -5654 -8190 -5650
rect -8186 -5654 -8168 -5650
rect -8164 -5654 -8138 -5650
rect -8134 -5654 -8116 -5650
rect -8112 -5654 -8086 -5650
rect -8082 -5654 -8064 -5650
rect -8060 -5654 -8057 -5650
rect -8245 -5656 -8057 -5654
rect -8034 -5654 -8030 -5648
rect -8002 -5654 -7998 -5648
rect -8235 -5662 -8231 -5656
rect -8183 -5662 -8179 -5656
rect -8131 -5662 -8127 -5656
rect -8079 -5662 -8075 -5656
rect -8258 -5711 -8235 -5706
rect -8258 -5777 -8253 -5711
rect -8227 -5715 -8223 -5702
rect -8235 -5719 -8223 -5715
rect -8205 -5711 -8183 -5706
rect -8235 -5724 -8231 -5719
rect -8240 -5773 -8235 -5768
rect -8227 -5777 -8223 -5764
rect -8205 -5777 -8200 -5711
rect -8175 -5715 -8171 -5702
rect -8123 -5706 -8119 -5702
rect -8071 -5706 -8067 -5702
rect -8026 -5706 -8022 -5694
rect -7994 -5706 -7990 -5694
rect -8183 -5719 -8171 -5715
rect -8153 -5711 -8131 -5706
rect -8123 -5711 -8079 -5706
rect -8071 -5711 -8034 -5706
rect -8026 -5711 -8002 -5706
rect -7994 -5711 -7946 -5706
rect -8183 -5724 -8179 -5719
rect -8188 -5773 -8183 -5768
rect -8175 -5777 -8171 -5764
rect -8153 -5777 -8148 -5711
rect -8134 -5734 -8131 -5729
rect -8123 -5738 -8119 -5711
rect -8131 -5769 -8127 -5758
rect -8131 -5773 -8119 -5769
rect -8258 -5782 -8235 -5777
rect -8227 -5782 -8183 -5777
rect -8175 -5782 -8131 -5777
rect -8227 -5785 -8223 -5782
rect -8175 -5785 -8171 -5782
rect -8123 -5785 -8119 -5773
rect -8101 -5777 -8096 -5711
rect -8082 -5734 -8079 -5729
rect -8071 -5738 -8067 -5711
rect -8026 -5714 -8022 -5711
rect -7994 -5714 -7990 -5711
rect -8034 -5741 -8030 -5734
rect -8002 -5741 -7998 -5734
rect -8044 -5743 -7980 -5741
rect -8044 -5747 -8042 -5743
rect -8038 -5747 -8018 -5743
rect -8014 -5747 -8010 -5743
rect -8006 -5747 -7986 -5743
rect -7982 -5747 -7980 -5743
rect -8044 -5749 -7980 -5747
rect -7951 -5748 -7946 -5711
rect -7929 -5718 -7924 -5462
rect -7898 -5443 -7892 -5442
rect -7898 -5447 -7897 -5443
rect -7893 -5447 -7892 -5443
rect -7898 -5450 -7892 -5447
rect -7863 -5450 -7858 -5439
rect -7813 -5445 -7804 -5442
rect -7813 -5449 -7811 -5445
rect -7807 -5449 -7804 -5445
rect -7813 -5450 -7804 -5449
rect -7898 -5454 -7886 -5450
rect -7898 -5464 -7892 -5454
rect -7828 -5454 -7804 -5450
rect -7750 -5446 -7746 -5438
rect -7697 -5444 -7643 -5441
rect -7863 -5462 -7848 -5458
rect -7813 -5462 -7804 -5454
rect -7778 -5458 -7765 -5454
rect -7778 -5461 -7774 -5458
rect -7898 -5468 -7897 -5464
rect -7893 -5468 -7892 -5464
rect -7898 -5469 -7892 -5468
rect -7863 -5472 -7858 -5462
rect -7813 -5466 -7811 -5462
rect -7807 -5466 -7804 -5462
rect -7813 -5469 -7804 -5466
rect -7786 -5472 -7782 -5469
rect -7834 -5476 -7782 -5472
rect -7834 -5481 -7830 -5476
rect -7892 -5486 -7830 -5481
rect -7898 -5494 -7892 -5493
rect -7898 -5498 -7897 -5494
rect -7893 -5498 -7892 -5494
rect -7898 -5501 -7892 -5498
rect -7863 -5501 -7858 -5486
rect -7778 -5492 -7774 -5469
rect -7771 -5476 -7765 -5458
rect -7697 -5448 -7694 -5444
rect -7690 -5448 -7677 -5444
rect -7673 -5448 -7667 -5444
rect -7663 -5448 -7650 -5444
rect -7646 -5448 -7643 -5444
rect -7697 -5450 -7643 -5448
rect -7742 -5476 -7738 -5466
rect -7689 -5475 -7685 -5450
rect -7654 -5475 -7650 -5450
rect -7771 -5481 -7750 -5476
rect -7742 -5481 -7724 -5476
rect -7742 -5484 -7738 -5481
rect -7813 -5496 -7804 -5493
rect -7813 -5500 -7811 -5496
rect -7807 -5500 -7804 -5496
rect -7813 -5501 -7804 -5500
rect -7898 -5505 -7886 -5501
rect -7898 -5515 -7892 -5505
rect -7828 -5505 -7804 -5501
rect -7863 -5513 -7848 -5509
rect -7813 -5513 -7804 -5505
rect -7898 -5519 -7897 -5515
rect -7893 -5519 -7892 -5515
rect -7898 -5520 -7892 -5519
rect -7863 -5524 -7858 -5513
rect -7813 -5517 -7811 -5513
rect -7807 -5517 -7804 -5513
rect -7813 -5520 -7804 -5517
rect -7786 -5524 -7782 -5502
rect -7750 -5504 -7746 -5494
rect -7729 -5501 -7724 -5481
rect -7758 -5505 -7731 -5504
rect -7758 -5509 -7757 -5505
rect -7753 -5509 -7736 -5505
rect -7732 -5509 -7731 -5505
rect -7758 -5510 -7731 -5509
rect -7728 -5518 -7724 -5501
rect -7863 -5527 -7782 -5524
rect -7729 -5538 -7724 -5518
rect -7702 -5517 -7689 -5512
rect -7681 -5515 -7677 -5495
rect -7662 -5515 -7658 -5495
rect -7650 -5511 -7643 -5507
rect -7702 -5522 -7697 -5517
rect -7681 -5519 -7658 -5515
rect -7648 -5519 -7643 -5511
rect -7635 -5514 -7608 -5511
rect -7635 -5518 -7632 -5514
rect -7628 -5518 -7615 -5514
rect -7611 -5518 -7608 -5514
rect -7702 -5527 -7671 -5522
rect -7702 -5538 -7697 -5527
rect -7729 -5543 -7706 -5538
rect -7701 -5543 -7697 -5538
rect -7662 -5539 -7658 -5519
rect -7635 -5520 -7608 -5518
rect -7627 -5525 -7623 -5520
rect -7866 -5624 -7812 -5621
rect -7866 -5628 -7863 -5624
rect -7859 -5628 -7846 -5624
rect -7842 -5628 -7836 -5624
rect -7832 -5628 -7819 -5624
rect -7815 -5628 -7812 -5624
rect -7866 -5630 -7812 -5628
rect -7858 -5655 -7854 -5630
rect -7823 -5655 -7819 -5630
rect -7871 -5697 -7858 -5692
rect -7850 -5695 -7846 -5675
rect -7831 -5695 -7827 -5675
rect -7819 -5691 -7812 -5687
rect -7871 -5702 -7866 -5697
rect -7850 -5699 -7827 -5695
rect -7817 -5699 -7812 -5691
rect -7804 -5694 -7777 -5691
rect -7804 -5698 -7801 -5694
rect -7797 -5698 -7784 -5694
rect -7780 -5698 -7777 -5694
rect -7871 -5707 -7840 -5702
rect -7871 -5718 -7866 -5707
rect -7929 -5723 -7866 -5718
rect -7831 -5719 -7827 -5699
rect -7804 -5700 -7777 -5698
rect -7796 -5705 -7792 -5700
rect -7831 -5725 -7808 -5719
rect -7831 -5729 -7827 -5725
rect -7951 -5753 -7911 -5748
rect -7839 -5755 -7835 -5749
rect -7814 -5755 -7808 -5725
rect -7729 -5738 -7724 -5543
rect -7662 -5545 -7639 -5539
rect -7662 -5549 -7658 -5545
rect -7670 -5575 -7666 -5569
rect -7645 -5575 -7639 -5545
rect -7619 -5575 -7615 -5565
rect -7670 -5579 -7658 -5575
rect -7697 -5601 -7684 -5596
rect -7678 -5601 -7672 -5596
rect -7697 -5734 -7692 -5601
rect -7662 -5604 -7658 -5579
rect -7645 -5580 -7627 -5575
rect -7619 -5580 -7588 -5575
rect -7619 -5592 -7615 -5580
rect -7627 -5609 -7623 -5603
rect -7635 -5610 -7608 -5609
rect -7635 -5614 -7634 -5610
rect -7630 -5614 -7613 -5610
rect -7609 -5614 -7608 -5610
rect -7635 -5615 -7608 -5614
rect -7670 -5630 -7666 -5624
rect -7678 -5631 -7651 -5630
rect -7678 -5635 -7677 -5631
rect -7673 -5635 -7656 -5631
rect -7652 -5635 -7651 -5631
rect -7678 -5636 -7651 -5635
rect -7593 -5687 -7588 -5580
rect -7549 -5648 -7522 -5645
rect -7549 -5652 -7546 -5648
rect -7542 -5652 -7529 -5648
rect -7525 -5652 -7522 -5648
rect -7549 -5654 -7522 -5652
rect -7541 -5666 -7537 -5654
rect -7593 -5692 -7583 -5687
rect -7576 -5689 -7553 -5687
rect -7576 -5692 -7541 -5689
rect -7558 -5694 -7541 -5692
rect -7533 -5698 -7529 -5686
rect -7431 -5686 -7427 -5211
rect -6992 -5613 -6928 -5610
rect -6992 -5617 -6989 -5613
rect -6985 -5617 -6967 -5613
rect -6963 -5617 -6957 -5613
rect -6953 -5617 -6935 -5613
rect -6931 -5617 -6928 -5613
rect -7193 -5621 -7005 -5618
rect -6992 -5619 -6928 -5617
rect -7193 -5625 -7190 -5621
rect -7186 -5625 -7168 -5621
rect -7164 -5625 -7138 -5621
rect -7134 -5625 -7116 -5621
rect -7112 -5625 -7086 -5621
rect -7082 -5625 -7064 -5621
rect -7060 -5625 -7034 -5621
rect -7030 -5625 -7012 -5621
rect -7008 -5625 -7005 -5621
rect -7193 -5627 -7005 -5625
rect -6982 -5625 -6978 -5619
rect -6950 -5625 -6946 -5619
rect -7183 -5633 -7179 -5627
rect -7131 -5633 -7127 -5627
rect -7079 -5633 -7075 -5627
rect -7027 -5633 -7023 -5627
rect -7307 -5681 -7303 -5673
rect -7206 -5682 -7183 -5677
rect -7431 -5690 -7366 -5686
rect -7541 -5702 -7529 -5698
rect -7500 -5696 -7473 -5693
rect -7500 -5700 -7497 -5696
rect -7493 -5700 -7480 -5696
rect -7476 -5700 -7473 -5696
rect -7500 -5702 -7473 -5700
rect -7541 -5714 -7537 -5702
rect -7492 -5710 -7488 -5702
rect -7370 -5706 -7366 -5690
rect -7370 -5709 -7314 -5706
rect -7370 -5710 -7306 -5709
rect -7587 -5739 -7557 -5738
rect -7587 -5743 -7556 -5739
rect -7788 -5755 -7784 -5745
rect -7587 -5755 -7582 -5743
rect -7565 -5744 -7556 -5743
rect -7533 -5740 -7529 -5733
rect -7484 -5740 -7480 -5730
rect -7317 -5713 -7306 -5710
rect -7317 -5723 -7314 -5713
rect -7299 -5714 -7295 -5701
rect -7317 -5736 -7314 -5728
rect -7307 -5729 -7303 -5724
rect -7289 -5729 -7288 -5725
rect -7206 -5735 -7201 -5682
rect -7175 -5686 -7171 -5673
rect -7183 -5690 -7171 -5686
rect -7153 -5682 -7131 -5677
rect -7183 -5695 -7179 -5690
rect -7317 -5740 -7307 -5736
rect -7533 -5745 -7492 -5740
rect -7484 -5745 -7421 -5740
rect -7228 -5741 -7201 -5735
rect -7533 -5748 -7529 -5745
rect -7484 -5748 -7480 -5745
rect -8079 -5769 -8075 -5758
rect -7839 -5759 -7827 -5755
rect -8079 -5773 -8067 -5769
rect -8101 -5782 -8079 -5777
rect -8071 -5785 -8067 -5773
rect -7866 -5776 -7860 -5774
rect -7866 -5781 -7853 -5776
rect -7847 -5781 -7841 -5776
rect -7831 -5784 -7827 -5759
rect -7814 -5760 -7796 -5755
rect -7788 -5760 -7608 -5755
rect -7602 -5760 -7582 -5755
rect -7548 -5752 -7511 -5748
rect -7548 -5758 -7544 -5752
rect -7515 -5758 -7511 -5752
rect -7788 -5772 -7784 -5760
rect -7492 -5768 -7488 -5758
rect -7796 -5789 -7792 -5783
rect -7556 -5775 -7552 -5768
rect -7523 -5775 -7519 -5768
rect -7500 -5769 -7473 -5768
rect -7500 -5773 -7499 -5769
rect -7495 -5773 -7478 -5769
rect -7474 -5773 -7473 -5769
rect -7500 -5774 -7473 -5773
rect -7564 -5776 -7537 -5775
rect -7564 -5780 -7563 -5776
rect -7559 -5780 -7542 -5776
rect -7538 -5780 -7537 -5776
rect -7564 -5781 -7537 -5780
rect -7531 -5776 -7504 -5775
rect -7531 -5780 -7530 -5776
rect -7526 -5780 -7509 -5776
rect -7505 -5780 -7504 -5776
rect -7531 -5781 -7504 -5780
rect -7426 -5787 -7421 -5745
rect -7206 -5748 -7201 -5741
rect -7188 -5744 -7183 -5739
rect -7175 -5748 -7171 -5735
rect -7153 -5748 -7148 -5682
rect -7123 -5686 -7119 -5673
rect -7071 -5677 -7067 -5673
rect -7019 -5677 -7015 -5673
rect -6974 -5677 -6970 -5665
rect -6942 -5677 -6938 -5665
rect -6831 -5674 -6804 -5671
rect -7131 -5690 -7119 -5686
rect -7101 -5682 -7079 -5677
rect -7071 -5682 -7027 -5677
rect -7019 -5682 -6982 -5677
rect -6974 -5682 -6950 -5677
rect -6942 -5682 -6874 -5677
rect -6831 -5678 -6828 -5674
rect -6824 -5678 -6811 -5674
rect -6807 -5678 -6804 -5674
rect -6831 -5680 -6804 -5678
rect -7131 -5695 -7127 -5690
rect -7136 -5744 -7131 -5739
rect -7123 -5748 -7119 -5735
rect -7101 -5748 -7096 -5682
rect -7082 -5705 -7079 -5700
rect -7071 -5709 -7067 -5682
rect -7079 -5740 -7075 -5729
rect -7079 -5744 -7067 -5740
rect -7299 -5757 -7295 -5756
rect -7324 -5760 -7295 -5757
rect -7299 -5763 -7295 -5760
rect -7289 -5763 -7285 -5756
rect -7328 -5767 -7306 -5763
rect -7299 -5767 -7285 -5763
rect -7328 -5768 -7311 -5767
rect -7328 -5787 -7323 -5768
rect -7804 -5790 -7777 -5789
rect -7804 -5794 -7803 -5790
rect -7799 -5794 -7782 -5790
rect -7778 -5794 -7777 -5790
rect -7804 -5795 -7777 -5794
rect -8235 -5813 -8231 -5805
rect -8183 -5813 -8179 -5805
rect -8131 -5813 -8127 -5805
rect -8079 -5813 -8075 -5805
rect -7839 -5810 -7835 -5804
rect -7847 -5811 -7820 -5810
rect -8245 -5814 -8057 -5813
rect -8245 -5818 -8218 -5814
rect -8214 -5818 -8166 -5814
rect -8162 -5818 -8114 -5814
rect -8110 -5818 -8062 -5814
rect -8058 -5818 -8057 -5814
rect -7847 -5815 -7846 -5811
rect -7842 -5815 -7825 -5811
rect -7821 -5815 -7820 -5811
rect -7847 -5816 -7820 -5815
rect -8245 -5819 -8057 -5818
rect -8252 -5832 -8245 -5827
rect -8240 -5832 -8193 -5827
rect -8188 -5832 -8139 -5827
rect -8134 -5832 -8087 -5827
rect -7697 -5838 -7692 -5789
rect -7635 -5797 -7631 -5787
rect -7426 -5792 -7323 -5787
rect -7314 -5787 -7311 -5768
rect -7299 -5768 -7295 -5767
rect -7289 -5768 -7285 -5767
rect -7206 -5753 -7183 -5748
rect -7175 -5753 -7131 -5748
rect -7123 -5753 -7079 -5748
rect -7175 -5756 -7171 -5753
rect -7123 -5756 -7119 -5753
rect -7071 -5756 -7067 -5744
rect -7049 -5748 -7044 -5682
rect -7030 -5705 -7027 -5700
rect -7019 -5709 -7015 -5682
rect -6974 -5685 -6970 -5682
rect -6942 -5685 -6938 -5682
rect -6982 -5712 -6978 -5705
rect -6950 -5712 -6946 -5705
rect -6992 -5714 -6928 -5712
rect -6992 -5718 -6990 -5714
rect -6986 -5718 -6966 -5714
rect -6962 -5718 -6958 -5714
rect -6954 -5718 -6934 -5714
rect -6930 -5718 -6928 -5714
rect -6992 -5720 -6928 -5718
rect -7027 -5740 -7023 -5729
rect -6879 -5736 -6874 -5682
rect -6823 -5685 -6819 -5680
rect -6815 -5735 -6811 -5725
rect -6833 -5736 -6823 -5735
rect -6879 -5740 -6823 -5736
rect -6815 -5740 -6802 -5735
rect -7027 -5744 -7015 -5740
rect -6879 -5741 -6829 -5740
rect -7049 -5753 -7027 -5748
rect -7019 -5756 -7015 -5744
rect -6815 -5752 -6811 -5740
rect -7281 -5763 -7277 -5756
rect -7281 -5767 -7265 -5763
rect -7281 -5768 -7277 -5767
rect -7307 -5779 -7303 -5778
rect -7290 -5783 -7282 -5779
rect -7278 -5783 -7276 -5779
rect -7268 -5787 -7265 -5767
rect -6823 -5769 -6819 -5763
rect -6831 -5770 -6804 -5769
rect -6831 -5774 -6830 -5770
rect -6826 -5774 -6809 -5770
rect -6805 -5774 -6804 -5770
rect -6831 -5775 -6804 -5774
rect -7183 -5784 -7179 -5776
rect -7131 -5784 -7127 -5776
rect -7079 -5784 -7075 -5776
rect -7027 -5784 -7023 -5776
rect -7314 -5790 -7265 -5787
rect -7193 -5785 -7005 -5784
rect -7193 -5789 -7166 -5785
rect -7162 -5789 -7114 -5785
rect -7110 -5789 -7062 -5785
rect -7058 -5789 -7010 -5785
rect -7006 -5789 -7005 -5785
rect -7193 -5790 -7005 -5789
rect -7200 -5803 -7193 -5798
rect -7188 -5803 -7141 -5798
rect -7136 -5803 -7087 -5798
rect -7082 -5803 -7035 -5798
rect -7645 -5829 -7634 -5825
rect -7715 -5843 -7692 -5838
rect -7661 -5834 -7642 -5829
rect -7627 -5830 -7623 -5817
rect -7661 -5843 -7656 -5834
rect -7715 -5924 -7710 -5843
rect -7697 -5848 -7656 -5843
rect -7645 -5839 -7642 -5834
rect -7645 -5852 -7642 -5844
rect -7635 -5845 -7631 -5840
rect -7617 -5845 -7616 -5841
rect -7645 -5856 -7635 -5852
rect -7269 -5853 -7205 -5850
rect -7269 -5857 -7266 -5853
rect -7262 -5857 -7244 -5853
rect -7240 -5857 -7234 -5853
rect -7230 -5857 -7212 -5853
rect -7208 -5857 -7205 -5853
rect -7470 -5861 -7282 -5858
rect -7269 -5859 -7205 -5857
rect -7470 -5865 -7467 -5861
rect -7463 -5865 -7445 -5861
rect -7441 -5865 -7415 -5861
rect -7411 -5865 -7393 -5861
rect -7389 -5865 -7363 -5861
rect -7359 -5865 -7341 -5861
rect -7337 -5865 -7311 -5861
rect -7307 -5865 -7289 -5861
rect -7285 -5865 -7282 -5861
rect -7470 -5867 -7282 -5865
rect -7259 -5865 -7255 -5859
rect -7227 -5865 -7223 -5859
rect -7627 -5878 -7623 -5872
rect -7617 -5878 -7613 -5872
rect -7654 -5911 -7648 -5882
rect -7642 -5883 -7634 -5879
rect -7627 -5883 -7613 -5878
rect -7642 -5886 -7639 -5883
rect -7627 -5884 -7623 -5883
rect -7617 -5884 -7613 -5883
rect -7609 -5879 -7605 -5872
rect -7460 -5873 -7456 -5867
rect -7408 -5873 -7404 -5867
rect -7356 -5873 -7352 -5867
rect -7304 -5873 -7300 -5867
rect -7609 -5883 -7593 -5879
rect -7609 -5884 -7605 -5883
rect -7642 -5903 -7639 -5891
rect -7635 -5895 -7631 -5894
rect -7618 -5899 -7610 -5895
rect -7606 -5899 -7604 -5895
rect -7596 -5903 -7593 -5883
rect -7642 -5906 -7593 -5903
rect -7654 -5917 -7478 -5911
rect -7132 -5896 -7105 -5893
rect -7132 -5900 -7129 -5896
rect -7125 -5900 -7112 -5896
rect -7108 -5900 -7105 -5896
rect -7132 -5902 -7105 -5900
rect -7484 -5922 -7460 -5917
rect -7715 -5929 -7570 -5924
rect -7669 -5953 -7605 -5950
rect -7669 -5957 -7666 -5953
rect -7662 -5957 -7644 -5953
rect -7640 -5957 -7634 -5953
rect -7630 -5957 -7612 -5953
rect -7608 -5957 -7605 -5953
rect -7870 -5961 -7682 -5958
rect -7669 -5959 -7605 -5957
rect -7870 -5965 -7867 -5961
rect -7863 -5965 -7845 -5961
rect -7841 -5965 -7815 -5961
rect -7811 -5965 -7793 -5961
rect -7789 -5965 -7763 -5961
rect -7759 -5965 -7741 -5961
rect -7737 -5965 -7711 -5961
rect -7707 -5965 -7689 -5961
rect -7685 -5965 -7682 -5961
rect -7870 -5967 -7682 -5965
rect -7659 -5965 -7655 -5959
rect -7627 -5965 -7623 -5959
rect -7860 -5973 -7856 -5967
rect -7808 -5973 -7804 -5967
rect -7756 -5973 -7752 -5967
rect -7704 -5973 -7700 -5967
rect -7883 -6022 -7860 -6017
rect -7883 -6088 -7878 -6022
rect -7852 -6026 -7848 -6013
rect -7860 -6030 -7848 -6026
rect -7830 -6022 -7808 -6017
rect -7860 -6035 -7856 -6030
rect -7865 -6084 -7860 -6079
rect -7852 -6088 -7848 -6075
rect -7830 -6088 -7825 -6022
rect -7800 -6026 -7796 -6013
rect -7748 -6017 -7744 -6013
rect -7696 -6017 -7692 -6013
rect -7651 -6017 -7647 -6005
rect -7619 -6017 -7615 -6005
rect -7575 -6017 -7570 -5929
rect -7484 -5931 -7478 -5922
rect -7452 -5926 -7448 -5913
rect -7483 -5988 -7478 -5931
rect -7460 -5930 -7448 -5926
rect -7430 -5922 -7408 -5917
rect -7460 -5935 -7456 -5930
rect -7465 -5984 -7460 -5979
rect -7452 -5988 -7448 -5975
rect -7430 -5988 -7425 -5922
rect -7400 -5926 -7396 -5913
rect -7348 -5917 -7344 -5913
rect -7296 -5917 -7292 -5913
rect -7251 -5917 -7247 -5905
rect -7219 -5917 -7215 -5905
rect -7124 -5907 -7120 -5902
rect -7408 -5930 -7396 -5926
rect -7378 -5922 -7356 -5917
rect -7348 -5922 -7304 -5917
rect -7296 -5922 -7259 -5917
rect -7251 -5922 -7227 -5917
rect -7219 -5922 -7162 -5917
rect -7408 -5935 -7404 -5930
rect -7413 -5984 -7408 -5979
rect -7400 -5988 -7396 -5975
rect -7378 -5988 -7373 -5922
rect -7359 -5945 -7356 -5940
rect -7348 -5949 -7344 -5922
rect -7356 -5980 -7352 -5969
rect -7356 -5984 -7344 -5980
rect -7483 -5993 -7460 -5988
rect -7452 -5993 -7408 -5988
rect -7400 -5993 -7356 -5988
rect -7452 -5996 -7448 -5993
rect -7400 -5996 -7396 -5993
rect -7348 -5996 -7344 -5984
rect -7326 -5988 -7321 -5922
rect -7307 -5945 -7304 -5940
rect -7296 -5949 -7292 -5922
rect -7251 -5925 -7247 -5922
rect -7219 -5925 -7215 -5922
rect -7259 -5952 -7255 -5945
rect -7227 -5952 -7223 -5945
rect -7269 -5954 -7205 -5952
rect -7269 -5958 -7267 -5954
rect -7263 -5958 -7243 -5954
rect -7239 -5958 -7235 -5954
rect -7231 -5958 -7211 -5954
rect -7207 -5958 -7205 -5954
rect -7269 -5960 -7205 -5958
rect -7167 -5958 -7162 -5922
rect -7116 -5957 -7112 -5947
rect -7134 -5958 -7124 -5957
rect -7167 -5962 -7124 -5958
rect -7116 -5962 -7103 -5957
rect -7167 -5963 -7131 -5962
rect -7304 -5980 -7300 -5969
rect -7116 -5974 -7112 -5962
rect -7304 -5984 -7292 -5980
rect -7326 -5993 -7304 -5988
rect -7296 -5996 -7292 -5984
rect -7124 -5991 -7120 -5985
rect -7808 -6030 -7796 -6026
rect -7778 -6022 -7756 -6017
rect -7748 -6022 -7704 -6017
rect -7696 -6022 -7659 -6017
rect -7651 -6022 -7627 -6017
rect -7619 -6022 -7570 -6017
rect -7132 -5992 -7105 -5991
rect -7132 -5996 -7131 -5992
rect -7127 -5996 -7110 -5992
rect -7106 -5996 -7105 -5992
rect -7132 -5997 -7105 -5996
rect -7808 -6035 -7804 -6030
rect -7813 -6084 -7808 -6079
rect -7800 -6088 -7796 -6075
rect -7778 -6088 -7773 -6022
rect -7759 -6045 -7756 -6040
rect -7748 -6049 -7744 -6022
rect -7756 -6080 -7752 -6069
rect -7756 -6084 -7744 -6080
rect -7883 -6093 -7860 -6088
rect -7852 -6093 -7808 -6088
rect -7800 -6093 -7756 -6088
rect -7852 -6096 -7848 -6093
rect -7800 -6096 -7796 -6093
rect -7748 -6096 -7744 -6084
rect -7726 -6088 -7721 -6022
rect -7707 -6045 -7704 -6040
rect -7696 -6049 -7692 -6022
rect -7651 -6025 -7647 -6022
rect -7619 -6025 -7615 -6022
rect -7659 -6052 -7655 -6045
rect -7627 -6052 -7623 -6045
rect -7669 -6054 -7605 -6052
rect -7669 -6058 -7667 -6054
rect -7663 -6058 -7643 -6054
rect -7639 -6058 -7635 -6054
rect -7631 -6058 -7611 -6054
rect -7607 -6058 -7605 -6054
rect -7669 -6060 -7605 -6058
rect -7704 -6080 -7700 -6069
rect -7704 -6084 -7692 -6080
rect -7726 -6093 -7704 -6088
rect -7696 -6096 -7692 -6084
rect -7860 -6124 -7856 -6116
rect -7808 -6124 -7804 -6116
rect -7756 -6124 -7752 -6116
rect -7704 -6124 -7700 -6116
rect -7870 -6125 -7682 -6124
rect -7870 -6129 -7843 -6125
rect -7839 -6129 -7791 -6125
rect -7787 -6129 -7739 -6125
rect -7735 -6129 -7687 -6125
rect -7683 -6129 -7682 -6125
rect -7870 -6130 -7682 -6129
rect -7877 -6143 -7870 -6138
rect -7865 -6143 -7818 -6138
rect -7813 -6143 -7764 -6138
rect -7759 -6143 -7712 -6138
rect -7577 -6205 -7572 -6022
rect -7460 -6024 -7456 -6016
rect -7408 -6024 -7404 -6016
rect -7356 -6024 -7352 -6016
rect -7304 -6024 -7300 -6016
rect -7470 -6025 -7282 -6024
rect -7470 -6029 -7443 -6025
rect -7439 -6029 -7391 -6025
rect -7387 -6029 -7339 -6025
rect -7335 -6029 -7287 -6025
rect -7283 -6029 -7282 -6025
rect -7470 -6030 -7282 -6029
rect -7477 -6043 -7470 -6038
rect -7465 -6043 -7418 -6038
rect -7413 -6043 -7364 -6038
rect -7359 -6043 -7312 -6038
rect -7556 -6141 -7529 -6138
rect -7556 -6145 -7553 -6141
rect -7549 -6145 -7536 -6141
rect -7532 -6145 -7529 -6141
rect -7556 -6147 -7529 -6145
rect -7548 -6152 -7544 -6147
rect -7540 -6202 -7536 -6192
rect -7558 -6205 -7548 -6202
rect -7577 -6207 -7548 -6205
rect -7540 -6207 -7527 -6202
rect -7577 -6210 -7555 -6207
rect -7540 -6219 -7536 -6207
rect -7548 -6236 -7544 -6230
rect -7556 -6237 -7529 -6236
rect -7556 -6241 -7555 -6237
rect -7551 -6241 -7534 -6237
rect -7530 -6241 -7529 -6237
rect -7556 -6242 -7529 -6241
<< m2contact >>
rect -2883 -554 -2877 -549
rect -2913 -636 -2907 -631
rect -2000 -779 -1995 -774
rect -1948 -779 -1943 -774
rect -1894 -740 -1889 -735
rect -1842 -740 -1837 -735
rect -2000 -838 -1995 -833
rect -1948 -838 -1943 -833
rect -1894 -838 -1889 -833
rect -1842 -838 -1837 -833
rect -8323 -3102 -8318 -3097
rect -7668 -3030 -7659 -3025
rect -8271 -3102 -8266 -3097
rect -8217 -3063 -8212 -3058
rect -8165 -3063 -8160 -3058
rect -8323 -3161 -8318 -3156
rect -8271 -3161 -8266 -3156
rect -8217 -3161 -8212 -3156
rect -8165 -3161 -8160 -3156
rect -8309 -3406 -8304 -3401
rect -7882 -3105 -7873 -3100
rect -7595 -3151 -7589 -3146
rect -7813 -3312 -7807 -3307
rect -8029 -3344 -8024 -3339
rect -8257 -3406 -8252 -3401
rect -8203 -3367 -8198 -3362
rect -8151 -3367 -8146 -3362
rect -7856 -3378 -7850 -3373
rect -7843 -3394 -7837 -3389
rect -7771 -3373 -7765 -3368
rect -8309 -3465 -8304 -3460
rect -8257 -3465 -8252 -3460
rect -8203 -3465 -8198 -3460
rect -8151 -3465 -8146 -3460
rect -7625 -3233 -7619 -3228
rect -7450 -3189 -7444 -3184
rect -7257 -3205 -7251 -3200
rect -7480 -3271 -7474 -3266
rect -7408 -3250 -7402 -3245
rect -7111 -3203 -7105 -3198
rect -6967 -3207 -6961 -3202
rect -7023 -3233 -7015 -3228
rect -7300 -3287 -7292 -3281
rect -7287 -3287 -7281 -3282
rect -7141 -3285 -7135 -3280
rect -6812 -3209 -6806 -3204
rect -7029 -3320 -7024 -3315
rect -6997 -3289 -6991 -3284
rect -6677 -3217 -6671 -3212
rect -6842 -3291 -6836 -3286
rect -6568 -3244 -6562 -3239
rect -6720 -3299 -6714 -3294
rect -6707 -3299 -6701 -3294
rect -6575 -3295 -6568 -3290
rect -6272 -3333 -6267 -3328
rect -6256 -3405 -6251 -3400
rect -6089 -3482 -6083 -3477
rect -5923 -3556 -5918 -3551
rect -5871 -3556 -5866 -3551
rect -5817 -3517 -5812 -3512
rect -5765 -3517 -5760 -3512
rect -5923 -3615 -5918 -3610
rect -5871 -3615 -5866 -3610
rect -5817 -3615 -5812 -3610
rect -5765 -3615 -5760 -3610
rect -7360 -3871 -7355 -3866
rect -7071 -3765 -7066 -3760
rect -8254 -4014 -8249 -4009
rect -8202 -4014 -8197 -4009
rect -8148 -3975 -8143 -3970
rect -8096 -3975 -8091 -3970
rect -8254 -4073 -8249 -4068
rect -8202 -4073 -8197 -4068
rect -8148 -4073 -8143 -4068
rect -8096 -4073 -8091 -4068
rect -8237 -4255 -8232 -4250
rect -8185 -4255 -8180 -4250
rect -8131 -4216 -8126 -4211
rect -8079 -4216 -8074 -4211
rect -7876 -3956 -7871 -3951
rect -7820 -4227 -7814 -4222
rect -7890 -4279 -7885 -4274
rect -7587 -3966 -7581 -3961
rect -7647 -3991 -7635 -3986
rect -7360 -3901 -7355 -3896
rect -7418 -3965 -7412 -3960
rect -7466 -3989 -7461 -3983
rect -7254 -3963 -7248 -3958
rect -7114 -3965 -7108 -3960
rect -7174 -3989 -7169 -3984
rect -7630 -4048 -7621 -4042
rect -7617 -4048 -7611 -4043
rect -7448 -4047 -7442 -4042
rect -7284 -4045 -7278 -4040
rect -6963 -3978 -6957 -3973
rect -7154 -4048 -7148 -4042
rect -7144 -4047 -7138 -4042
rect -7048 -4026 -7041 -4021
rect -6993 -4060 -6987 -4055
rect -6718 -4041 -6708 -4036
rect -6800 -4182 -6794 -4177
rect -7241 -4259 -7236 -4254
rect -6866 -4257 -6861 -4252
rect -6830 -4264 -6824 -4259
rect -7863 -4292 -7857 -4287
rect -7850 -4309 -7844 -4304
rect -8237 -4314 -8232 -4309
rect -8185 -4314 -8180 -4309
rect -8131 -4314 -8126 -4309
rect -8079 -4314 -8074 -4309
rect -6450 -4411 -6443 -4406
rect -6185 -4378 -6180 -4373
rect -6218 -4427 -6212 -4421
rect -6198 -4449 -6193 -4444
rect -6185 -4449 -6180 -4444
rect -6166 -4449 -6161 -4444
rect -6144 -4477 -6138 -4471
rect -6090 -4481 -6085 -4476
rect -6038 -4481 -6033 -4476
rect -5984 -4442 -5979 -4437
rect -5932 -4442 -5927 -4437
rect -6090 -4540 -6085 -4535
rect -6038 -4540 -6033 -4535
rect -5984 -4540 -5979 -4535
rect -5932 -4540 -5927 -4535
rect -8248 -4818 -8243 -4813
rect -7876 -4724 -7871 -4719
rect -8196 -4818 -8191 -4813
rect -8142 -4779 -8137 -4774
rect -8090 -4779 -8085 -4774
rect -8248 -4877 -8243 -4872
rect -8196 -4877 -8191 -4872
rect -8142 -4877 -8137 -4872
rect -8090 -4877 -8085 -4872
rect -8235 -5130 -8230 -5125
rect -7976 -5068 -7970 -5063
rect -8183 -5130 -8178 -5125
rect -8129 -5091 -8124 -5086
rect -8077 -5091 -8072 -5086
rect -7826 -5076 -7820 -5071
rect -7566 -4739 -7560 -4734
rect -7637 -4764 -7632 -4759
rect -7628 -4764 -7623 -4759
rect -7660 -4805 -7651 -4798
rect -7596 -4821 -7590 -4816
rect -7565 -4944 -7559 -4939
rect -7621 -4968 -7616 -4963
rect -7608 -5026 -7602 -5021
rect -7595 -5026 -7589 -5021
rect -7331 -5015 -7321 -5010
rect -7125 -4990 -7120 -4985
rect -7103 -4989 -7098 -4984
rect -7690 -5119 -7685 -5114
rect -7134 -5037 -7129 -5032
rect -7116 -5060 -7111 -5055
rect -7103 -5060 -7098 -5055
rect -7084 -5060 -7079 -5055
rect -7067 -5094 -7062 -5089
rect -7009 -5090 -7004 -5085
rect -6957 -5090 -6952 -5085
rect -6903 -5051 -6898 -5046
rect -6851 -5051 -6846 -5046
rect -3978 -5089 -3973 -5084
rect -7869 -5143 -7863 -5138
rect -7856 -5158 -7850 -5153
rect -7690 -5153 -7685 -5148
rect -7009 -5149 -7004 -5144
rect -6957 -5149 -6952 -5144
rect -6903 -5149 -6898 -5144
rect -6851 -5149 -6846 -5144
rect -8235 -5189 -8230 -5184
rect -8183 -5189 -8178 -5184
rect -8129 -5189 -8124 -5184
rect -8077 -5189 -8072 -5184
rect -3991 -5160 -3986 -5155
rect -3978 -5160 -3973 -5155
rect -3959 -5160 -3954 -5155
rect -7661 -5302 -7652 -5295
rect -7584 -5302 -7576 -5295
rect -8248 -5524 -8243 -5519
rect -8196 -5524 -8191 -5519
rect -8142 -5485 -8137 -5480
rect -8090 -5485 -8085 -5480
rect -8248 -5583 -8243 -5578
rect -8196 -5583 -8191 -5578
rect -8142 -5583 -8137 -5578
rect -8090 -5583 -8085 -5578
rect -8245 -5773 -8240 -5768
rect -8193 -5773 -8188 -5768
rect -8139 -5734 -8134 -5729
rect -8087 -5734 -8082 -5729
rect -7898 -5486 -7892 -5481
rect -7654 -5519 -7648 -5514
rect -7706 -5543 -7701 -5538
rect -7823 -5699 -7817 -5694
rect -7911 -5753 -7906 -5748
rect -7729 -5743 -7724 -5738
rect -7684 -5601 -7678 -5596
rect -7583 -5692 -7576 -5687
rect -7697 -5744 -7692 -5734
rect -7295 -5713 -7290 -5708
rect -7234 -5741 -7228 -5735
rect -7866 -5774 -7860 -5769
rect -7853 -5781 -7847 -5776
rect -7608 -5760 -7602 -5755
rect -7697 -5789 -7692 -5774
rect -7193 -5744 -7188 -5739
rect -7141 -5744 -7136 -5739
rect -7087 -5705 -7082 -5700
rect -7324 -5757 -7319 -5751
rect -8245 -5832 -8240 -5827
rect -8193 -5832 -8188 -5827
rect -8139 -5832 -8134 -5827
rect -8087 -5832 -8082 -5827
rect -7035 -5705 -7030 -5700
rect -7308 -5784 -7303 -5779
rect -7295 -5784 -7290 -5779
rect -7276 -5784 -7271 -5779
rect -7193 -5803 -7188 -5798
rect -7141 -5803 -7136 -5798
rect -7087 -5803 -7082 -5798
rect -7035 -5803 -7030 -5798
rect -7623 -5829 -7618 -5824
rect -7654 -5882 -7648 -5877
rect -7644 -5891 -7639 -5886
rect -7636 -5900 -7631 -5895
rect -7623 -5900 -7618 -5895
rect -7604 -5900 -7599 -5895
rect -7870 -6084 -7865 -6079
rect -7470 -5984 -7465 -5979
rect -7418 -5984 -7413 -5979
rect -7364 -5945 -7359 -5940
rect -7312 -5945 -7307 -5940
rect -7818 -6084 -7813 -6079
rect -7764 -6045 -7759 -6040
rect -7712 -6045 -7707 -6040
rect -7870 -6143 -7865 -6138
rect -7818 -6143 -7813 -6138
rect -7764 -6143 -7759 -6138
rect -7712 -6143 -7707 -6138
rect -7470 -6043 -7465 -6038
rect -7418 -6043 -7413 -6038
rect -7364 -6043 -7359 -6038
rect -7312 -6043 -7307 -6038
<< metal2 >>
rect -2883 -619 -2877 -554
rect -2913 -626 -2877 -619
rect -2913 -631 -2907 -626
rect -2000 -833 -1995 -779
rect -1948 -833 -1943 -779
rect -1894 -833 -1889 -740
rect -1842 -833 -1837 -740
rect -7691 -2963 -6122 -2958
rect -8323 -3156 -8318 -3102
rect -8271 -3156 -8266 -3102
rect -8217 -3156 -8212 -3063
rect -8165 -3156 -8160 -3063
rect -7896 -3105 -7882 -3100
rect -7896 -3106 -7873 -3105
rect -8024 -3344 -7999 -3339
rect -8309 -3460 -8304 -3406
rect -8257 -3460 -8252 -3406
rect -8203 -3460 -8198 -3367
rect -8151 -3460 -8146 -3367
rect -8004 -3373 -7999 -3344
rect -7896 -3373 -7890 -3106
rect -8004 -3379 -7856 -3373
rect -7813 -3377 -7807 -3312
rect -7691 -3368 -7686 -2963
rect -7668 -3035 -7659 -3030
rect -7765 -3373 -7686 -3368
rect -7843 -3384 -7807 -3377
rect -7843 -3389 -7837 -3384
rect -7664 -3760 -7659 -3035
rect -7395 -3068 -6592 -3063
rect -7595 -3216 -7589 -3151
rect -7625 -3223 -7589 -3216
rect -7625 -3228 -7619 -3223
rect -7450 -3254 -7444 -3189
rect -7395 -3245 -7390 -3068
rect -6751 -3098 -6611 -3093
rect -7402 -3250 -7390 -3245
rect -7480 -3261 -7444 -3254
rect -7480 -3266 -7474 -3261
rect -7257 -3270 -7251 -3205
rect -7111 -3268 -7105 -3203
rect -7287 -3277 -7251 -3270
rect -7141 -3275 -7105 -3268
rect -7041 -3233 -7023 -3228
rect -7353 -3287 -7300 -3281
rect -7287 -3282 -7281 -3277
rect -7141 -3280 -7135 -3275
rect -7353 -3288 -7292 -3287
rect -7353 -3675 -7346 -3288
rect -7041 -3360 -7036 -3233
rect -6967 -3272 -6961 -3207
rect -6997 -3279 -6961 -3272
rect -6812 -3274 -6806 -3209
rect -6997 -3284 -6991 -3279
rect -6842 -3281 -6806 -3274
rect -6842 -3286 -6836 -3281
rect -7029 -3346 -7024 -3320
rect -6751 -3346 -6746 -3098
rect -6677 -3282 -6671 -3217
rect -6707 -3289 -6671 -3282
rect -7029 -3351 -6746 -3346
rect -6734 -3294 -6714 -3293
rect -6734 -3299 -6720 -3294
rect -6707 -3294 -6701 -3289
rect -6616 -3290 -6611 -3098
rect -6597 -3239 -6592 -3068
rect -6597 -3244 -6568 -3239
rect -6616 -3295 -6575 -3290
rect -6734 -3300 -6714 -3299
rect -7041 -3365 -6890 -3360
rect -7353 -3682 -7041 -3675
rect -7664 -3765 -7071 -3760
rect -7485 -3862 -7169 -3857
rect -7890 -3956 -7876 -3951
rect -8254 -4068 -8249 -4014
rect -8202 -4068 -8197 -4014
rect -8148 -4068 -8143 -3975
rect -8096 -4068 -8091 -3975
rect -8237 -4309 -8232 -4255
rect -8185 -4309 -8180 -4255
rect -8131 -4309 -8126 -4216
rect -8079 -4309 -8074 -4216
rect -7890 -4274 -7885 -3956
rect -7647 -4025 -7643 -3991
rect -7650 -4027 -7643 -4025
rect -7650 -4029 -7644 -4027
rect -7719 -4035 -7644 -4029
rect -7587 -4031 -7581 -3966
rect -7485 -3996 -7480 -3862
rect -7360 -3896 -7355 -3871
rect -7466 -3996 -7461 -3989
rect -7485 -4001 -7461 -3996
rect -7890 -4287 -7885 -4279
rect -7890 -4292 -7863 -4287
rect -7820 -4292 -7814 -4227
rect -7850 -4299 -7814 -4292
rect -7850 -4304 -7844 -4299
rect -7889 -4724 -7876 -4719
rect -8248 -4872 -8243 -4818
rect -8196 -4872 -8191 -4818
rect -8142 -4872 -8137 -4779
rect -8090 -4872 -8085 -4779
rect -7970 -5068 -7959 -5063
rect -8235 -5184 -8230 -5130
rect -8183 -5184 -8178 -5130
rect -8129 -5184 -8124 -5091
rect -8077 -5184 -8072 -5091
rect -7964 -5113 -7959 -5068
rect -7889 -5113 -7884 -4724
rect -7964 -5118 -7884 -5113
rect -7889 -5138 -7884 -5118
rect -7889 -5143 -7869 -5138
rect -7826 -5141 -7820 -5076
rect -7856 -5148 -7820 -5141
rect -7856 -5153 -7850 -5148
rect -8248 -5578 -8243 -5524
rect -8196 -5578 -8191 -5524
rect -8142 -5578 -8137 -5485
rect -8090 -5578 -8085 -5485
rect -7911 -5486 -7898 -5481
rect -8245 -5827 -8240 -5773
rect -8193 -5827 -8188 -5773
rect -8139 -5827 -8134 -5734
rect -8087 -5827 -8082 -5734
rect -7911 -5748 -7906 -5486
rect -7911 -5769 -7906 -5753
rect -7823 -5764 -7817 -5699
rect -7911 -5774 -7866 -5769
rect -7853 -5771 -7817 -5764
rect -7853 -5776 -7847 -5771
rect -7729 -5891 -7724 -5743
rect -7719 -5747 -7713 -4035
rect -7617 -4038 -7581 -4031
rect -7647 -4048 -7630 -4042
rect -7617 -4043 -7611 -4038
rect -7647 -4049 -7639 -4048
rect -7709 -4805 -7660 -4798
rect -7709 -5295 -7703 -4805
rect -7690 -5148 -7685 -5119
rect -7709 -5302 -7661 -5295
rect -7647 -5393 -7643 -4049
rect -7466 -4632 -7461 -4001
rect -7418 -4030 -7412 -3965
rect -7254 -4028 -7248 -3963
rect -7174 -3984 -7169 -3862
rect -7448 -4037 -7412 -4030
rect -7284 -4035 -7248 -4028
rect -7114 -4030 -7108 -3965
rect -7048 -4021 -7041 -3682
rect -7448 -4042 -7442 -4037
rect -7284 -4040 -7278 -4035
rect -7144 -4037 -7108 -4030
rect -7144 -4042 -7138 -4037
rect -6963 -4043 -6957 -3978
rect -7154 -4093 -7148 -4048
rect -6993 -4050 -6957 -4043
rect -6993 -4055 -6987 -4050
rect -6895 -4054 -6890 -3365
rect -6734 -3550 -6727 -3300
rect -6272 -3400 -6267 -3333
rect -6272 -3405 -6256 -3400
rect -6127 -3477 -6122 -2963
rect -6127 -3482 -6089 -3477
rect -6734 -3557 -6700 -3550
rect -6707 -3848 -6700 -3557
rect -5923 -3610 -5918 -3556
rect -5871 -3610 -5866 -3556
rect -5817 -3610 -5812 -3517
rect -5765 -3610 -5760 -3517
rect -6707 -3855 -6443 -3848
rect -6901 -4059 -6890 -4054
rect -6866 -4036 -6713 -4033
rect -6866 -4038 -6718 -4036
rect -7628 -4637 -7461 -4632
rect -7454 -4099 -7148 -4093
rect -7628 -4759 -7623 -4637
rect -7454 -4647 -7448 -4099
rect -6901 -4199 -6896 -4059
rect -7503 -4653 -7448 -4647
rect -7327 -4204 -6896 -4199
rect -7637 -4963 -7632 -4764
rect -7566 -4804 -7560 -4739
rect -7596 -4811 -7560 -4804
rect -7596 -4816 -7590 -4811
rect -7637 -4968 -7621 -4963
rect -7565 -5009 -7559 -4944
rect -7595 -5016 -7559 -5009
rect -7595 -5021 -7589 -5016
rect -7706 -5397 -7643 -5393
rect -7608 -5078 -7602 -5026
rect -7503 -5078 -7497 -4653
rect -7327 -5010 -7322 -4204
rect -6866 -4252 -6861 -4038
rect -6725 -4041 -6718 -4038
rect -6800 -4247 -6794 -4182
rect -6866 -4258 -6861 -4257
rect -6830 -4254 -6794 -4247
rect -7241 -4832 -7236 -4259
rect -6830 -4259 -6824 -4254
rect -6450 -4406 -6443 -3855
rect -6180 -4377 -6162 -4374
rect -6218 -4471 -6212 -4427
rect -6165 -4444 -6162 -4377
rect -6193 -4448 -6185 -4444
rect -6218 -4477 -6144 -4471
rect -6090 -4535 -6085 -4481
rect -6038 -4535 -6033 -4481
rect -5984 -4535 -5979 -4442
rect -5932 -4535 -5927 -4442
rect -7241 -4837 -7182 -4832
rect -7187 -4962 -7182 -4837
rect -7187 -4967 -7144 -4962
rect -7149 -4985 -7144 -4967
rect -7149 -4990 -7125 -4985
rect -7098 -4988 -7080 -4985
rect -7608 -5084 -7497 -5078
rect -7706 -5538 -7702 -5397
rect -7654 -5584 -7648 -5519
rect -7684 -5591 -7648 -5584
rect -7684 -5596 -7678 -5591
rect -7697 -5747 -7692 -5744
rect -7719 -5752 -7692 -5747
rect -7697 -5774 -7692 -5752
rect -7608 -5755 -7602 -5084
rect -7134 -5089 -7129 -5037
rect -7083 -5055 -7080 -4988
rect -7111 -5059 -7103 -5055
rect -7134 -5094 -7067 -5089
rect -7009 -5144 -7004 -5090
rect -6957 -5144 -6952 -5090
rect -6903 -5144 -6898 -5051
rect -6851 -5144 -6846 -5051
rect -3973 -5088 -3955 -5085
rect -3958 -5155 -3955 -5088
rect -3986 -5159 -3978 -5155
rect -7583 -5687 -7576 -5302
rect -7290 -5712 -7272 -5709
rect -7608 -5761 -7602 -5760
rect -7351 -5757 -7324 -5751
rect -7351 -5809 -7345 -5757
rect -7275 -5779 -7272 -5712
rect -7303 -5783 -7295 -5779
rect -7234 -5809 -7228 -5741
rect -7193 -5798 -7188 -5744
rect -7141 -5798 -7136 -5744
rect -7087 -5798 -7082 -5705
rect -7035 -5798 -7030 -5705
rect -7351 -5815 -7228 -5809
rect -7618 -5828 -7600 -5825
rect -7648 -5882 -7617 -5878
rect -7635 -5883 -7617 -5882
rect -7675 -5891 -7644 -5886
rect -7729 -5896 -7670 -5891
rect -7603 -5895 -7600 -5828
rect -7631 -5899 -7623 -5895
rect -7470 -6038 -7465 -5984
rect -7870 -6138 -7865 -6084
rect -7818 -6138 -7813 -6084
rect -7764 -6138 -7759 -6045
rect -7418 -6038 -7413 -5984
rect -7364 -6038 -7359 -5945
rect -7312 -6038 -7307 -5945
rect -7712 -6138 -7707 -6045
<< m123contact >>
rect -6207 -4393 -6202 -4388
rect -6184 -4394 -6179 -4389
rect -7125 -5004 -7120 -4999
rect -7102 -5005 -7097 -5000
rect -4000 -5104 -3995 -5099
rect -3977 -5105 -3972 -5100
rect -7317 -5728 -7312 -5723
rect -7294 -5729 -7289 -5724
rect -7645 -5844 -7640 -5839
rect -7622 -5845 -7617 -5840
<< metal3 >>
rect -6202 -4393 -6184 -4389
rect -7120 -5004 -7102 -5000
rect -3995 -5104 -3977 -5100
rect -7312 -5728 -7294 -5724
rect -7640 -5844 -7622 -5840
<< labels >>
rlabel metal1 -2587 -601 -2587 -601 3 gnd
rlabel metal1 -2501 -601 -2501 -601 7 vdd
rlabel metal1 -2501 -652 -2501 -652 7 vdd
rlabel metal1 -2587 -652 -2587 -652 3 gnd
rlabel metal1 -2437 -580 -2437 -580 5 vdd
rlabel metal1 -2437 -653 -2437 -653 1 gnd
rlabel metal1 -2234 -763 -2234 -763 1 gnd
rlabel metal1 -2234 -690 -2234 -690 5 vdd
rlabel metal1 -2283 -642 -2283 -642 5 vdd
rlabel metal1 -2298 -770 -2298 -770 1 gnd
rlabel metal1 -2265 -770 -2265 -770 1 gnd
rlabel metal1 -2851 -647 -2851 -647 1 gnd
rlabel metal1 -2851 -551 -2851 -551 5 vdd
rlabel metal1 -2886 -481 -2886 -481 5 vdd
rlabel metal1 -2913 -481 -2913 -481 5 vdd
rlabel metal1 -2894 -668 -2894 -668 1 gnd
rlabel metal1 -7895 -5455 -7895 -5455 3 gnd
rlabel metal1 -7809 -5455 -7809 -5455 7 vdd
rlabel metal1 -7809 -5506 -7809 -5506 7 vdd
rlabel metal1 -7895 -5506 -7895 -5506 3 gnd
rlabel metal1 -7745 -5434 -7745 -5434 5 vdd
rlabel metal1 -7745 -5507 -7745 -5507 1 gnd
rlabel metal1 -7873 -4693 -7873 -4693 3 gnd
rlabel metal1 -7787 -4693 -7787 -4693 7 vdd
rlabel metal1 -7787 -4744 -7787 -4744 7 vdd
rlabel metal1 -7873 -4744 -7873 -4744 3 gnd
rlabel metal1 -7723 -4672 -7723 -4672 5 vdd
rlabel metal1 -7723 -4745 -7723 -4745 1 gnd
rlabel metal1 -7873 -3925 -7873 -3925 3 gnd
rlabel metal1 -7787 -3925 -7787 -3925 7 vdd
rlabel metal1 -7787 -3976 -7787 -3976 7 vdd
rlabel metal1 -7873 -3976 -7873 -3976 3 gnd
rlabel metal1 -7723 -3904 -7723 -3904 5 vdd
rlabel metal1 -7723 -3977 -7723 -3977 1 gnd
rlabel metal1 -7879 -3074 -7879 -3074 3 gnd
rlabel metal1 -7793 -3074 -7793 -3074 7 vdd
rlabel metal1 -7793 -3125 -7793 -3125 7 vdd
rlabel metal1 -7879 -3125 -7879 -3125 3 gnd
rlabel metal1 -7729 -3053 -7729 -3053 5 vdd
rlabel metal1 -7729 -3126 -7729 -3126 1 gnd
rlabel metal1 -7831 -4341 -7831 -4341 1 gnd
rlabel metal1 -7850 -4154 -7850 -4154 5 vdd
rlabel metal1 -7823 -4154 -7823 -4154 5 vdd
rlabel metal1 -7788 -4224 -7788 -4224 5 vdd
rlabel metal1 -7788 -4320 -7788 -4320 1 gnd
rlabel metal1 -7837 -5190 -7837 -5190 1 gnd
rlabel metal1 -7856 -5003 -7856 -5003 5 vdd
rlabel metal1 -7829 -5003 -7829 -5003 5 vdd
rlabel metal1 -7794 -5073 -7794 -5073 5 vdd
rlabel metal1 -7794 -5169 -7794 -5169 1 gnd
rlabel metal1 -7715 -3097 -7715 -3097 1 p3
rlabel metal1 -7781 -3405 -7781 -3405 1 gnd
rlabel metal1 -7781 -3309 -7781 -3309 5 vdd
rlabel metal1 -7816 -3239 -7816 -3239 5 vdd
rlabel metal1 -7843 -3239 -7843 -3239 5 vdd
rlabel metal1 -7824 -3426 -7824 -3426 1 gnd
rlabel metal1 -7834 -5813 -7834 -5813 1 gnd
rlabel metal1 -7853 -5626 -7853 -5626 5 vdd
rlabel metal1 -7826 -5626 -7826 -5626 5 vdd
rlabel metal1 -7791 -5696 -7791 -5696 5 vdd
rlabel metal1 -7791 -5792 -7791 -5792 1 gnd
rlabel metal1 -7731 -5478 -7731 -5478 1 p0
rlabel metal1 -7779 -5757 -7779 -5757 1 g0
rlabel metal1 -7665 -5633 -7665 -5633 1 gnd
rlabel metal1 -7684 -5446 -7684 -5446 5 vdd
rlabel metal1 -7657 -5446 -7657 -5446 5 vdd
rlabel metal1 -7622 -5516 -7622 -5516 5 vdd
rlabel metal1 -7622 -5612 -7622 -5612 1 gnd
rlabel metal1 -7518 -5778 -7518 -5778 1 gnd
rlabel metal1 -7551 -5778 -7551 -5778 1 gnd
rlabel metal1 -7536 -5650 -7536 -5650 5 vdd
rlabel metal1 -7487 -5698 -7487 -5698 5 vdd
rlabel metal1 -7487 -5771 -7487 -5771 1 gnd
rlabel metal1 -7474 -5742 -7474 -5742 1 c1
rlabel metal1 -7577 -4853 -7577 -4853 1 gnd
rlabel metal1 -7596 -4666 -7596 -4666 5 vdd
rlabel metal1 -7569 -4666 -7569 -4666 5 vdd
rlabel metal1 -7534 -4736 -7534 -4736 5 vdd
rlabel metal1 -7534 -4832 -7534 -4832 1 gnd
rlabel metal1 -7576 -5058 -7576 -5058 1 gnd
rlabel metal1 -7595 -4871 -7595 -4871 5 vdd
rlabel metal1 -7568 -4871 -7568 -4871 5 vdd
rlabel metal1 -7533 -4941 -7533 -4941 5 vdd
rlabel metal1 -7533 -5037 -7533 -5037 1 gnd
rlabel metal1 -7782 -5134 -7782 -5134 1 g1
rlabel metal1 -7521 -4797 -7521 -4797 1 0c2
rlabel metal1 -7519 -5003 -7519 -5003 1 1c2
rlabel metal1 -7381 -4928 -7381 -4928 1 gnd
rlabel metal1 -7381 -4855 -7381 -4855 5 vdd
rlabel metal1 -7430 -4807 -7430 -4807 5 vdd
rlabel metal1 -7445 -4935 -7445 -4935 1 gnd
rlabel metal1 -7412 -4935 -7412 -4935 1 gnd
rlabel metal1 -7235 -5041 -7235 -5041 1 gnd
rlabel metal1 -7235 -4968 -7235 -4968 5 vdd
rlabel metal1 -7284 -4920 -7284 -4920 5 vdd
rlabel metal1 -7299 -5048 -7299 -5048 1 gnd
rlabel metal1 -7266 -5048 -7266 -5048 1 gnd
rlabel metal1 -7343 -4900 -7343 -4900 1 2c2
rlabel metal1 -7221 -5012 -7221 -5012 1 c2
rlabel metal1 -7555 -4059 -7555 -4059 1 gnd
rlabel metal1 -7555 -3963 -7555 -3963 5 vdd
rlabel metal1 -7590 -3893 -7590 -3893 5 vdd
rlabel metal1 -7617 -3893 -7617 -3893 5 vdd
rlabel metal1 -7598 -4080 -7598 -4080 1 gnd
rlabel metal1 -7429 -4079 -7429 -4079 1 gnd
rlabel metal1 -7448 -3892 -7448 -3892 5 vdd
rlabel metal1 -7421 -3892 -7421 -3892 5 vdd
rlabel metal1 -7386 -3962 -7386 -3962 5 vdd
rlabel metal1 -7386 -4058 -7386 -4058 1 gnd
rlabel metal1 -7265 -4077 -7265 -4077 1 gnd
rlabel metal1 -7284 -3890 -7284 -3890 5 vdd
rlabel metal1 -7257 -3890 -7257 -3890 5 vdd
rlabel metal1 -7222 -3960 -7222 -3960 5 vdd
rlabel metal1 -7222 -4056 -7222 -4056 1 gnd
rlabel metal1 -7710 -3949 -7710 -3949 1 p2
rlabel metal1 -7774 -4286 -7774 -4286 1 g2
rlabel metal1 -7525 -4024 -7525 -4024 1 0c3
rlabel metal1 -7372 -4024 -7372 -4024 1 1c3
rlabel metal1 -7208 -4021 -7208 -4021 1 2c3
rlabel metal1 -7082 -4058 -7082 -4058 1 gnd
rlabel metal1 -7082 -3962 -7082 -3962 5 vdd
rlabel metal1 -7117 -3892 -7117 -3892 5 vdd
rlabel metal1 -7144 -3892 -7144 -3892 5 vdd
rlabel metal1 -7125 -4079 -7125 -4079 1 gnd
rlabel metal1 -6768 -4275 -6768 -4275 1 gnd
rlabel metal1 -6768 -4179 -6768 -4179 5 vdd
rlabel metal1 -6803 -4109 -6803 -4109 5 vdd
rlabel metal1 -6830 -4109 -6830 -4109 5 vdd
rlabel metal1 -6811 -4296 -6811 -4296 1 gnd
rlabel metal1 -7067 -4024 -7067 -4024 1 3c3
rlabel metal1 -6754 -4241 -6754 -4241 1 5c3
rlabel metal1 -6665 -4075 -6665 -4075 1 gnd
rlabel metal1 -6698 -4075 -6698 -4075 1 gnd
rlabel metal1 -6683 -3947 -6683 -3947 5 vdd
rlabel metal1 -6634 -3995 -6634 -3995 5 vdd
rlabel metal1 -6634 -4068 -6634 -4068 1 gnd
rlabel metal1 -6500 -4278 -6500 -4278 1 gnd
rlabel metal1 -6500 -4205 -6500 -4205 5 vdd
rlabel metal1 -6549 -4157 -6549 -4157 5 vdd
rlabel metal1 -6564 -4285 -6564 -4285 1 gnd
rlabel metal1 -6531 -4285 -6531 -4285 1 gnd
rlabel metal1 -6353 -4438 -6353 -4438 1 gnd
rlabel metal1 -6353 -4365 -6353 -4365 5 vdd
rlabel metal1 -6402 -4317 -6402 -4317 5 vdd
rlabel metal1 -6417 -4445 -6417 -4445 1 gnd
rlabel metal1 -6384 -4445 -6384 -4445 1 gnd
rlabel metal1 -6622 -4039 -6622 -4039 1 6c3
rlabel metal1 -6485 -4250 -6485 -4250 1 7c3
rlabel metal1 -6339 -4409 -6339 -4409 1 c3
rlabel metal1 -7563 -3244 -7563 -3244 1 gnd
rlabel metal1 -7563 -3148 -7563 -3148 5 vdd
rlabel metal1 -7598 -3078 -7598 -3078 5 vdd
rlabel metal1 -7625 -3078 -7625 -3078 5 vdd
rlabel metal1 -7606 -3265 -7606 -3265 1 gnd
rlabel metal1 -7550 -3209 -7550 -3209 1 2c4
rlabel metal1 -7461 -3303 -7461 -3303 1 gnd
rlabel metal1 -7480 -3116 -7480 -3116 5 vdd
rlabel metal1 -7453 -3116 -7453 -3116 5 vdd
rlabel metal1 -7418 -3186 -7418 -3186 5 vdd
rlabel metal1 -7418 -3282 -7418 -3282 1 gnd
rlabel m2contact -7404 -3248 -7404 -3248 1 3c3
rlabel metal1 -7225 -3298 -7225 -3298 1 gnd
rlabel metal1 -7225 -3202 -7225 -3202 5 vdd
rlabel metal1 -7260 -3132 -7260 -3132 5 vdd
rlabel metal1 -7287 -3132 -7287 -3132 5 vdd
rlabel metal1 -7268 -3319 -7268 -3319 1 gnd
rlabel metal1 -7079 -3296 -7079 -3296 1 gnd
rlabel metal1 -7079 -3200 -7079 -3200 5 vdd
rlabel metal1 -7114 -3130 -7114 -3130 5 vdd
rlabel metal1 -7141 -3130 -7141 -3130 5 vdd
rlabel metal1 -7122 -3317 -7122 -3317 1 gnd
rlabel metal1 -7212 -3263 -7212 -3263 1 5c4
rlabel metal1 -7065 -3261 -7065 -3261 1 6c4
rlabel metal1 -6935 -3300 -6935 -3300 1 gnd
rlabel metal1 -6935 -3204 -6935 -3204 5 vdd
rlabel metal1 -6970 -3134 -6970 -3134 5 vdd
rlabel metal1 -6997 -3134 -6997 -3134 5 vdd
rlabel metal1 -6978 -3321 -6978 -3321 1 gnd
rlabel metal1 -6780 -3302 -6780 -3302 1 gnd
rlabel metal1 -6780 -3206 -6780 -3206 5 vdd
rlabel metal1 -6815 -3136 -6815 -3136 5 vdd
rlabel metal1 -6842 -3136 -6842 -3136 5 vdd
rlabel metal1 -6823 -3323 -6823 -3323 1 gnd
rlabel metal1 -6931 -4071 -6931 -4071 1 gnd
rlabel metal1 -6931 -3975 -6931 -3975 5 vdd
rlabel metal1 -6966 -3905 -6966 -3905 5 vdd
rlabel metal1 -6993 -3905 -6993 -3905 5 vdd
rlabel metal1 -6974 -4092 -6974 -4092 1 gnd
rlabel metal1 -6918 -4037 -6918 -4037 1 4c3
rlabel metal1 -6921 -3265 -6921 -3265 1 7c4
rlabel metal1 -6766 -3268 -6766 -3268 1 8c4
rlabel metal1 -6645 -3310 -6645 -3310 1 gnd
rlabel metal1 -6645 -3214 -6645 -3214 5 vdd
rlabel metal1 -6680 -3144 -6680 -3144 5 vdd
rlabel metal1 -6707 -3144 -6707 -3144 5 vdd
rlabel metal1 -6688 -3331 -6688 -3331 1 gnd
rlabel metal1 -6631 -3275 -6631 -3275 1 9c4
rlabel metal1 -6497 -3321 -6497 -3321 1 gnd
rlabel metal1 -6497 -3248 -6497 -3248 5 vdd
rlabel metal1 -6546 -3200 -6546 -3200 5 vdd
rlabel metal1 -6561 -3328 -6561 -3328 1 gnd
rlabel metal1 -6528 -3328 -6528 -3328 1 gnd
rlabel metal1 -6366 -3384 -6366 -3384 1 gnd
rlabel metal1 -6399 -3384 -6399 -3384 1 gnd
rlabel metal1 -6384 -3256 -6384 -3256 5 vdd
rlabel metal1 -6335 -3304 -6335 -3304 5 vdd
rlabel metal1 -6335 -3377 -6335 -3377 1 gnd
rlabel metal1 -6208 -3440 -6208 -3440 1 gnd
rlabel metal1 -6241 -3440 -6241 -3440 1 gnd
rlabel metal1 -6226 -3312 -6226 -3312 5 vdd
rlabel metal1 -6177 -3360 -6177 -3360 5 vdd
rlabel metal1 -6177 -3433 -6177 -3433 1 gnd
rlabel metal1 -6042 -3516 -6042 -3516 1 gnd
rlabel metal1 -6075 -3516 -6075 -3516 1 gnd
rlabel metal1 -6060 -3388 -6060 -3388 5 vdd
rlabel metal1 -6011 -3436 -6011 -3436 5 vdd
rlabel metal1 -6011 -3509 -6011 -3509 1 gnd
rlabel metal1 -6483 -3293 -6483 -3293 1 10c4
rlabel metal1 -6322 -3348 -6322 -3348 1 11c4
rlabel metal1 -6164 -3405 -6164 -3405 1 12c4
rlabel m2contact -7767 -3370 -7767 -3370 1 g3
rlabel metal1 -3995 -5088 -3993 -5086 3 a
rlabel metal1 -3995 -5142 -3993 -5140 1 b
rlabel metal1 -3989 -5105 -3987 -5104 1 gnd
rlabel metal1 -3989 -5050 -3987 -5048 5 vdd
rlabel metal1 -3977 -5142 -3973 -5140 1 out
rlabel metal1 -3981 -5088 -3979 -5085 1 a_bar
rlabel metal1 -7306 -5729 -7304 -5728 1 gnd
rlabel metal1 -7298 -5712 -7296 -5709 1 a_bar
rlabel metal1 -7414 -5688 -7414 -5688 1 p1
rlabel metal1 -7634 -5845 -7632 -5844 1 gnd
rlabel metal1 -7634 -5790 -7632 -5788 5 vdd
rlabel metal1 -7626 -5828 -7624 -5825 1 a_bar
rlabel metal1 -7114 -5005 -7112 -5004 1 gnd
rlabel metal1 -7114 -4950 -7112 -4948 5 vdd
rlabel metal1 -7106 -4988 -7104 -4985 1 a_bar
rlabel metal1 -6196 -4394 -6194 -4393 1 gnd
rlabel metal1 -6196 -4339 -6194 -4337 5 vdd
rlabel metal1 -6188 -4377 -6186 -4374 1 a_bar
rlabel metal1 -8018 -5460 -8018 -5460 1 qnot
rlabel metal1 -8053 -5460 -8053 -5460 1 qmid
rlabel metal1 -8072 -5529 -8072 -5529 1 d4
rlabel metal1 -8101 -5493 -8101 -5493 1 b
rlabel metal1 -8124 -5528 -8124 -5528 1 d3
rlabel metal1 -8154 -5492 -8154 -5492 1 q1
rlabel metal1 -8176 -5460 -8176 -5460 1 d2
rlabel metal1 -8206 -5491 -8206 -5491 1 a
rlabel metal1 -8228 -5461 -8228 -5461 1 d1
rlabel metal1 -8253 -5581 -8253 -5581 1 clk
rlabel metal1 -8031 -5394 -8031 -5394 5 vdd
rlabel metal1 -8032 -5496 -8032 -5496 1 gnd
rlabel metal1 -7999 -5394 -7999 -5394 5 vdd
rlabel metal1 -8000 -5496 -8000 -5496 1 gnd
rlabel metal1 -8076 -5402 -8076 -5402 5 vdd
rlabel metal1 -8076 -5567 -8076 -5567 1 gnd
rlabel metal1 -8128 -5402 -8128 -5402 5 vdd
rlabel metal1 -8128 -5567 -8128 -5567 1 gnd
rlabel metal1 -8180 -5567 -8180 -5567 1 gnd
rlabel metal1 -8180 -5402 -8180 -5402 5 vdd
rlabel metal1 -8232 -5567 -8232 -5567 1 gnd
rlabel metal1 -8232 -5402 -8232 -5402 5 vdd
rlabel metal1 -8229 -5651 -8229 -5651 5 vdd
rlabel metal1 -8229 -5816 -8229 -5816 1 gnd
rlabel metal1 -8177 -5651 -8177 -5651 5 vdd
rlabel metal1 -8177 -5816 -8177 -5816 1 gnd
rlabel metal1 -8125 -5816 -8125 -5816 1 gnd
rlabel metal1 -8125 -5651 -8125 -5651 5 vdd
rlabel metal1 -8073 -5816 -8073 -5816 1 gnd
rlabel metal1 -8073 -5651 -8073 -5651 5 vdd
rlabel metal1 -7997 -5745 -7997 -5745 1 gnd
rlabel metal1 -7996 -5643 -7996 -5643 5 vdd
rlabel metal1 -8029 -5745 -8029 -5745 1 gnd
rlabel metal1 -8028 -5643 -8028 -5643 5 vdd
rlabel metal1 -8250 -5830 -8250 -5830 1 clk
rlabel metal1 -8225 -5710 -8225 -5710 1 d1
rlabel metal1 -8203 -5740 -8203 -5740 1 a
rlabel metal1 -8173 -5709 -8173 -5709 1 d2
rlabel metal1 -8151 -5741 -8151 -5741 1 q1
rlabel metal1 -8121 -5777 -8121 -5777 1 d3
rlabel metal1 -8098 -5742 -8098 -5742 1 b
rlabel metal1 -8069 -5778 -8069 -5778 1 d4
rlabel metal1 -8050 -5709 -8050 -5709 1 qmid
rlabel metal1 -8015 -5709 -8015 -5709 1 qnot
rlabel metal1 -8005 -5066 -8005 -5066 1 qnot
rlabel metal1 -8040 -5066 -8040 -5066 1 qmid
rlabel metal1 -8059 -5135 -8059 -5135 1 d4
rlabel metal1 -8088 -5099 -8088 -5099 1 b
rlabel metal1 -8111 -5134 -8111 -5134 1 d3
rlabel metal1 -8141 -5098 -8141 -5098 1 q1
rlabel metal1 -8163 -5066 -8163 -5066 1 d2
rlabel metal1 -8193 -5097 -8193 -5097 1 a
rlabel metal1 -8215 -5067 -8215 -5067 1 d1
rlabel metal1 -8240 -5187 -8240 -5187 1 clk
rlabel metal1 -8018 -5000 -8018 -5000 5 vdd
rlabel metal1 -8019 -5102 -8019 -5102 1 gnd
rlabel metal1 -7986 -5000 -7986 -5000 5 vdd
rlabel metal1 -7987 -5102 -7987 -5102 1 gnd
rlabel metal1 -8063 -5008 -8063 -5008 5 vdd
rlabel metal1 -8063 -5173 -8063 -5173 1 gnd
rlabel metal1 -8115 -5008 -8115 -5008 5 vdd
rlabel metal1 -8115 -5173 -8115 -5173 1 gnd
rlabel metal1 -8167 -5173 -8167 -5173 1 gnd
rlabel metal1 -8167 -5008 -8167 -5008 5 vdd
rlabel metal1 -8219 -5173 -8219 -5173 1 gnd
rlabel metal1 -8219 -5008 -8219 -5008 5 vdd
rlabel metal1 -8018 -4754 -8018 -4754 1 qnot
rlabel metal1 -8053 -4754 -8053 -4754 1 qmid
rlabel metal1 -8072 -4823 -8072 -4823 1 d4
rlabel metal1 -8101 -4787 -8101 -4787 1 b
rlabel metal1 -8124 -4822 -8124 -4822 1 d3
rlabel metal1 -8154 -4786 -8154 -4786 1 q1
rlabel metal1 -8176 -4754 -8176 -4754 1 d2
rlabel metal1 -8206 -4785 -8206 -4785 1 a
rlabel metal1 -8228 -4755 -8228 -4755 1 d1
rlabel metal1 -8253 -4875 -8253 -4875 1 clk
rlabel metal1 -8031 -4688 -8031 -4688 5 vdd
rlabel metal1 -8032 -4790 -8032 -4790 1 gnd
rlabel metal1 -7999 -4688 -7999 -4688 5 vdd
rlabel metal1 -8000 -4790 -8000 -4790 1 gnd
rlabel metal1 -8076 -4696 -8076 -4696 5 vdd
rlabel metal1 -8076 -4861 -8076 -4861 1 gnd
rlabel metal1 -8128 -4696 -8128 -4696 5 vdd
rlabel metal1 -8128 -4861 -8128 -4861 1 gnd
rlabel metal1 -8180 -4861 -8180 -4861 1 gnd
rlabel metal1 -8180 -4696 -8180 -4696 5 vdd
rlabel metal1 -8232 -4861 -8232 -4861 1 gnd
rlabel metal1 -8232 -4696 -8232 -4696 5 vdd
rlabel metal1 -8221 -4133 -8221 -4133 5 vdd
rlabel metal1 -8221 -4298 -8221 -4298 1 gnd
rlabel metal1 -8169 -4133 -8169 -4133 5 vdd
rlabel metal1 -8169 -4298 -8169 -4298 1 gnd
rlabel metal1 -8117 -4298 -8117 -4298 1 gnd
rlabel metal1 -8117 -4133 -8117 -4133 5 vdd
rlabel metal1 -8065 -4298 -8065 -4298 1 gnd
rlabel metal1 -8065 -4133 -8065 -4133 5 vdd
rlabel metal1 -7989 -4227 -7989 -4227 1 gnd
rlabel metal1 -7988 -4125 -7988 -4125 5 vdd
rlabel metal1 -8021 -4227 -8021 -4227 1 gnd
rlabel metal1 -8020 -4125 -8020 -4125 5 vdd
rlabel metal1 -8242 -4312 -8242 -4312 1 clk
rlabel metal1 -8217 -4192 -8217 -4192 1 d1
rlabel metal1 -8195 -4222 -8195 -4222 1 a
rlabel metal1 -8165 -4191 -8165 -4191 1 d2
rlabel metal1 -8143 -4223 -8143 -4223 1 q1
rlabel metal1 -8113 -4259 -8113 -4259 1 d3
rlabel metal1 -8090 -4224 -8090 -4224 1 b
rlabel metal1 -8061 -4260 -8061 -4260 1 d4
rlabel metal1 -8042 -4191 -8042 -4191 1 qmid
rlabel metal1 -8007 -4191 -8007 -4191 1 qnot
rlabel metal1 -8238 -3892 -8238 -3892 5 vdd
rlabel metal1 -8238 -4057 -8238 -4057 1 gnd
rlabel metal1 -8186 -3892 -8186 -3892 5 vdd
rlabel metal1 -8186 -4057 -8186 -4057 1 gnd
rlabel metal1 -8134 -4057 -8134 -4057 1 gnd
rlabel metal1 -8134 -3892 -8134 -3892 5 vdd
rlabel metal1 -8082 -4057 -8082 -4057 1 gnd
rlabel metal1 -8082 -3892 -8082 -3892 5 vdd
rlabel metal1 -8006 -3986 -8006 -3986 1 gnd
rlabel metal1 -8005 -3884 -8005 -3884 5 vdd
rlabel metal1 -8038 -3986 -8038 -3986 1 gnd
rlabel metal1 -8037 -3884 -8037 -3884 5 vdd
rlabel metal1 -8259 -4071 -8259 -4071 1 clk
rlabel metal1 -8234 -3951 -8234 -3951 1 d1
rlabel metal1 -8212 -3981 -8212 -3981 1 a
rlabel metal1 -8182 -3950 -8182 -3950 1 d2
rlabel metal1 -8160 -3982 -8160 -3982 1 q1
rlabel metal1 -8130 -4018 -8130 -4018 1 d3
rlabel metal1 -8107 -3983 -8107 -3983 1 b
rlabel metal1 -8078 -4019 -8078 -4019 1 d4
rlabel metal1 -8059 -3950 -8059 -3950 1 qmid
rlabel metal1 -8024 -3950 -8024 -3950 1 qnot
rlabel metal1 -8307 -2980 -8307 -2980 5 vdd
rlabel metal1 -8307 -3145 -8307 -3145 1 gnd
rlabel metal1 -8255 -2980 -8255 -2980 5 vdd
rlabel metal1 -8255 -3145 -8255 -3145 1 gnd
rlabel metal1 -8203 -3145 -8203 -3145 1 gnd
rlabel metal1 -8203 -2980 -8203 -2980 5 vdd
rlabel metal1 -8151 -3145 -8151 -3145 1 gnd
rlabel metal1 -8151 -2980 -8151 -2980 5 vdd
rlabel metal1 -8075 -3074 -8075 -3074 1 gnd
rlabel metal1 -8074 -2972 -8074 -2972 5 vdd
rlabel metal1 -8107 -3074 -8107 -3074 1 gnd
rlabel metal1 -8106 -2972 -8106 -2972 5 vdd
rlabel metal1 -8328 -3159 -8328 -3159 1 clk
rlabel metal1 -8303 -3039 -8303 -3039 1 d1
rlabel metal1 -8281 -3069 -8281 -3069 1 a
rlabel metal1 -8251 -3038 -8251 -3038 1 d2
rlabel metal1 -8229 -3070 -8229 -3070 1 q1
rlabel metal1 -8199 -3106 -8199 -3106 1 d3
rlabel metal1 -8176 -3071 -8176 -3071 1 b
rlabel metal1 -8147 -3107 -8147 -3107 1 d4
rlabel metal1 -8128 -3038 -8128 -3038 1 qmid
rlabel metal1 -8093 -3038 -8093 -3038 1 qnot
rlabel metal1 -8293 -3284 -8293 -3284 5 vdd
rlabel metal1 -8293 -3449 -8293 -3449 1 gnd
rlabel metal1 -8241 -3284 -8241 -3284 5 vdd
rlabel metal1 -8241 -3449 -8241 -3449 1 gnd
rlabel metal1 -8189 -3449 -8189 -3449 1 gnd
rlabel metal1 -8189 -3284 -8189 -3284 5 vdd
rlabel metal1 -8137 -3449 -8137 -3449 1 gnd
rlabel metal1 -8137 -3284 -8137 -3284 5 vdd
rlabel metal1 -8061 -3378 -8061 -3378 1 gnd
rlabel metal1 -8060 -3276 -8060 -3276 5 vdd
rlabel metal1 -8093 -3378 -8093 -3378 1 gnd
rlabel metal1 -8092 -3276 -8092 -3276 5 vdd
rlabel metal1 -8314 -3463 -8314 -3463 1 clk
rlabel metal1 -8289 -3343 -8289 -3343 1 d1
rlabel metal1 -8267 -3373 -8267 -3373 1 a
rlabel metal1 -8237 -3342 -8237 -3342 1 d2
rlabel metal1 -8215 -3374 -8215 -3374 1 q1
rlabel metal1 -8185 -3410 -8185 -3410 1 d3
rlabel metal1 -8162 -3375 -8162 -3375 1 b
rlabel metal1 -8133 -3411 -8133 -3411 1 d4
rlabel metal1 -8114 -3342 -8114 -3342 1 qmid
rlabel metal1 -8079 -3342 -8079 -3342 1 qnot
rlabel metal1 -7640 -6020 -7640 -6020 1 qnot
rlabel metal1 -7675 -6020 -7675 -6020 1 qmid
rlabel metal1 -7694 -6089 -7694 -6089 1 d4
rlabel metal1 -7723 -6053 -7723 -6053 1 b
rlabel metal1 -7746 -6088 -7746 -6088 1 d3
rlabel metal1 -7776 -6052 -7776 -6052 1 q1
rlabel metal1 -7798 -6020 -7798 -6020 1 d2
rlabel metal1 -7828 -6051 -7828 -6051 1 a
rlabel metal1 -7850 -6021 -7850 -6021 1 d1
rlabel metal1 -7875 -6141 -7875 -6141 1 clk
rlabel metal1 -7653 -5954 -7653 -5954 5 vdd
rlabel metal1 -7654 -6056 -7654 -6056 1 gnd
rlabel metal1 -7621 -5954 -7621 -5954 5 vdd
rlabel metal1 -7622 -6056 -7622 -6056 1 gnd
rlabel metal1 -7698 -5962 -7698 -5962 5 vdd
rlabel metal1 -7698 -6127 -7698 -6127 1 gnd
rlabel metal1 -7750 -5962 -7750 -5962 5 vdd
rlabel metal1 -7750 -6127 -7750 -6127 1 gnd
rlabel metal1 -7802 -6127 -7802 -6127 1 gnd
rlabel metal1 -7802 -5962 -7802 -5962 5 vdd
rlabel metal1 -7854 -6127 -7854 -6127 1 gnd
rlabel metal1 -7854 -5962 -7854 -5962 5 vdd
rlabel metal1 -7240 -5920 -7240 -5920 1 qnot
rlabel metal1 -7275 -5920 -7275 -5920 1 qmid
rlabel metal1 -7294 -5989 -7294 -5989 1 d4
rlabel metal1 -7323 -5953 -7323 -5953 1 b
rlabel metal1 -7346 -5988 -7346 -5988 1 d3
rlabel metal1 -7376 -5952 -7376 -5952 1 q1
rlabel metal1 -7398 -5920 -7398 -5920 1 d2
rlabel metal1 -7428 -5951 -7428 -5951 1 a
rlabel metal1 -7450 -5921 -7450 -5921 1 d1
rlabel metal1 -7475 -6041 -7475 -6041 1 clk
rlabel metal1 -7253 -5854 -7253 -5854 5 vdd
rlabel metal1 -7254 -5956 -7254 -5956 1 gnd
rlabel metal1 -7221 -5854 -7221 -5854 5 vdd
rlabel metal1 -7222 -5956 -7222 -5956 1 gnd
rlabel metal1 -7298 -5862 -7298 -5862 5 vdd
rlabel metal1 -7298 -6027 -7298 -6027 1 gnd
rlabel metal1 -7350 -5862 -7350 -5862 5 vdd
rlabel metal1 -7350 -6027 -7350 -6027 1 gnd
rlabel metal1 -7402 -6027 -7402 -6027 1 gnd
rlabel metal1 -7402 -5862 -7402 -5862 5 vdd
rlabel metal1 -7454 -6027 -7454 -6027 1 gnd
rlabel metal1 -7454 -5862 -7454 -5862 5 vdd
rlabel metal1 -6963 -5680 -6963 -5680 1 qnot
rlabel metal1 -6998 -5680 -6998 -5680 1 qmid
rlabel metal1 -7017 -5749 -7017 -5749 1 d4
rlabel metal1 -7046 -5713 -7046 -5713 1 b
rlabel metal1 -7069 -5748 -7069 -5748 1 d3
rlabel metal1 -7099 -5712 -7099 -5712 1 q1
rlabel metal1 -7121 -5680 -7121 -5680 1 d2
rlabel metal1 -7151 -5711 -7151 -5711 1 a
rlabel metal1 -7173 -5681 -7173 -5681 1 d1
rlabel metal1 -7198 -5801 -7198 -5801 1 clk
rlabel metal1 -6976 -5614 -6976 -5614 5 vdd
rlabel metal1 -6977 -5716 -6977 -5716 1 gnd
rlabel metal1 -6944 -5614 -6944 -5614 5 vdd
rlabel metal1 -6945 -5716 -6945 -5716 1 gnd
rlabel metal1 -7021 -5622 -7021 -5622 5 vdd
rlabel metal1 -7021 -5787 -7021 -5787 1 gnd
rlabel metal1 -7073 -5622 -7073 -5622 5 vdd
rlabel metal1 -7073 -5787 -7073 -5787 1 gnd
rlabel metal1 -7125 -5787 -7125 -5787 1 gnd
rlabel metal1 -7125 -5622 -7125 -5622 5 vdd
rlabel metal1 -7177 -5787 -7177 -5787 1 gnd
rlabel metal1 -7177 -5622 -7177 -5622 5 vdd
rlabel metal1 -6993 -4968 -6993 -4968 5 vdd
rlabel metal1 -6993 -5133 -6993 -5133 1 gnd
rlabel metal1 -6941 -4968 -6941 -4968 5 vdd
rlabel metal1 -6941 -5133 -6941 -5133 1 gnd
rlabel metal1 -6889 -5133 -6889 -5133 1 gnd
rlabel metal1 -6889 -4968 -6889 -4968 5 vdd
rlabel metal1 -6837 -5133 -6837 -5133 1 gnd
rlabel metal1 -6837 -4968 -6837 -4968 5 vdd
rlabel metal1 -6761 -5062 -6761 -5062 1 gnd
rlabel metal1 -6760 -4960 -6760 -4960 5 vdd
rlabel metal1 -6793 -5062 -6793 -5062 1 gnd
rlabel metal1 -6792 -4960 -6792 -4960 5 vdd
rlabel metal1 -7014 -5147 -7014 -5147 1 clk
rlabel metal1 -6989 -5027 -6989 -5027 1 d1
rlabel metal1 -6967 -5057 -6967 -5057 1 a
rlabel metal1 -6937 -5026 -6937 -5026 1 d2
rlabel metal1 -6915 -5058 -6915 -5058 1 q1
rlabel metal1 -6885 -5094 -6885 -5094 1 d3
rlabel metal1 -6862 -5059 -6862 -5059 1 b
rlabel metal1 -6833 -5095 -6833 -5095 1 d4
rlabel metal1 -6814 -5026 -6814 -5026 1 qmid
rlabel metal1 -6779 -5026 -6779 -5026 1 qnot
rlabel metal1 -6074 -4359 -6074 -4359 5 vdd
rlabel metal1 -6074 -4524 -6074 -4524 1 gnd
rlabel metal1 -6022 -4359 -6022 -4359 5 vdd
rlabel metal1 -6022 -4524 -6022 -4524 1 gnd
rlabel metal1 -5970 -4524 -5970 -4524 1 gnd
rlabel metal1 -5970 -4359 -5970 -4359 5 vdd
rlabel metal1 -5918 -4524 -5918 -4524 1 gnd
rlabel metal1 -5918 -4359 -5918 -4359 5 vdd
rlabel metal1 -5842 -4453 -5842 -4453 1 gnd
rlabel metal1 -5841 -4351 -5841 -4351 5 vdd
rlabel metal1 -5874 -4453 -5874 -4453 1 gnd
rlabel metal1 -5873 -4351 -5873 -4351 5 vdd
rlabel metal1 -6095 -4538 -6095 -4538 1 clk
rlabel metal1 -6070 -4418 -6070 -4418 1 d1
rlabel metal1 -6048 -4448 -6048 -4448 1 a
rlabel metal1 -6018 -4417 -6018 -4417 1 d2
rlabel metal1 -5996 -4449 -5996 -4449 1 q1
rlabel metal1 -5966 -4485 -5966 -4485 1 d3
rlabel metal1 -5943 -4450 -5943 -4450 1 b
rlabel metal1 -5914 -4486 -5914 -4486 1 d4
rlabel metal1 -5895 -4417 -5895 -4417 1 qmid
rlabel metal1 -5860 -4417 -5860 -4417 1 qnot
rlabel metal1 -5907 -3434 -5907 -3434 5 vdd
rlabel metal1 -5907 -3599 -5907 -3599 1 gnd
rlabel metal1 -5855 -3434 -5855 -3434 5 vdd
rlabel metal1 -5855 -3599 -5855 -3599 1 gnd
rlabel metal1 -5803 -3599 -5803 -3599 1 gnd
rlabel metal1 -5803 -3434 -5803 -3434 5 vdd
rlabel metal1 -5751 -3599 -5751 -3599 1 gnd
rlabel metal1 -5751 -3434 -5751 -3434 5 vdd
rlabel metal1 -5675 -3528 -5675 -3528 1 gnd
rlabel metal1 -5674 -3426 -5674 -3426 5 vdd
rlabel metal1 -5707 -3528 -5707 -3528 1 gnd
rlabel metal1 -5706 -3426 -5706 -3426 5 vdd
rlabel metal1 -5928 -3613 -5928 -3613 1 clk
rlabel metal1 -5903 -3493 -5903 -3493 1 d1
rlabel metal1 -5881 -3523 -5881 -3523 1 a
rlabel metal1 -5851 -3492 -5851 -3492 1 d2
rlabel metal1 -5829 -3524 -5829 -3524 1 q1
rlabel metal1 -5799 -3560 -5799 -3560 1 d3
rlabel metal1 -5776 -3525 -5776 -3525 1 b
rlabel metal1 -5747 -3561 -5747 -3561 1 d4
rlabel metal1 -5728 -3492 -5728 -3492 1 qmid
rlabel metal1 -5693 -3492 -5693 -3492 1 qnot
rlabel metal1 -7881 -6048 -7881 -6048 1 c0
rlabel metal1 -5660 -3492 -5660 -3492 1 c4
rlabel metal1 -8320 -3351 -8320 -3351 1 b3
rlabel metal1 -8334 -3054 -8334 -3054 3 a3
rlabel metal1 -8266 -3965 -8266 -3965 1 a2
rlabel metal1 -8248 -4213 -8248 -4213 1 b2
rlabel metal1 -8259 -4773 -8259 -4773 1 a1
rlabel metal1 -8246 -5093 -8246 -5093 1 b1
rlabel metal1 -8258 -5476 -8258 -5476 1 a0
rlabel metal1 -8256 -5738 -8256 -5738 1 b0
rlabel metal1 -7208 -5919 -7208 -5919 1 s0
rlabel metal1 -6929 -5679 -6929 -5679 1 s1
rlabel metal1 -6745 -5026 -6745 -5026 1 s2
rlabel metal1 -5827 -4416 -5827 -4416 1 s3
rlabel metal1 -1770 -715 -1770 -715 1 qnot
rlabel metal1 -1805 -715 -1805 -715 1 qmid
rlabel metal1 -1824 -784 -1824 -784 1 d4
rlabel metal1 -1853 -748 -1853 -748 1 b
rlabel metal1 -1876 -783 -1876 -783 1 d3
rlabel metal1 -1906 -747 -1906 -747 1 q1
rlabel metal1 -1928 -715 -1928 -715 1 d2
rlabel metal1 -1958 -746 -1958 -746 1 a
rlabel metal1 -1980 -716 -1980 -716 1 d1
rlabel metal1 -2005 -836 -2005 -836 1 clk
rlabel metal1 -1783 -649 -1783 -649 5 vdd
rlabel metal1 -1784 -751 -1784 -751 1 gnd
rlabel metal1 -1751 -649 -1751 -649 5 vdd
rlabel metal1 -1752 -751 -1752 -751 1 gnd
rlabel metal1 -1828 -657 -1828 -657 5 vdd
rlabel metal1 -1828 -822 -1828 -822 1 gnd
rlabel metal1 -1880 -657 -1880 -657 5 vdd
rlabel metal1 -1880 -822 -1880 -822 1 gnd
rlabel metal1 -1932 -822 -1932 -822 1 gnd
rlabel metal1 -1932 -657 -1932 -657 5 vdd
rlabel metal1 -1984 -822 -1984 -822 1 gnd
rlabel metal1 -1984 -657 -1984 -657 5 vdd
rlabel metal1 -5540 -3469 -5540 -3469 5 vdd
rlabel metal1 -5540 -3565 -5540 -3565 1 gnd
rlabel metal1 -5716 -4477 -5716 -4477 1 gnd
rlabel metal1 -5716 -4381 -5716 -4381 5 vdd
rlabel metal1 -6682 -5097 -6682 -5097 1 gnd
rlabel metal1 -6682 -5001 -6682 -5001 5 vdd
rlabel metal1 -6818 -5772 -6818 -5772 1 gnd
rlabel metal1 -6818 -5676 -6818 -5676 5 vdd
rlabel metal1 -7119 -5994 -7119 -5994 1 gnd
rlabel metal1 -7119 -5898 -7119 -5898 5 vdd
rlabel metal1 -7543 -6239 -7543 -6239 1 gnd
rlabel metal1 -7543 -6143 -7543 -6143 5 vdd
<< end >>
